module Ctrl(
  input        io_cacheCtrl_iCache_stall, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_fetchUnit_allow_to_go, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_decodeUnit_inst0_src1_ren, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input  [4:0] io_decodeUnit_inst0_src1_raddr, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_decodeUnit_inst0_src2_ren, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input  [4:0] io_decodeUnit_inst0_src2_raddr, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_decodeUnit_branch, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_decodeUnit_allow_to_go, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_decodeUnit_do_flush, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_executeUnit_inst_0_is_load, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input  [4:0] io_executeUnit_inst_0_reg_waddr, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_executeUnit_inst_1_is_load, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input  [4:0] io_executeUnit_inst_1_reg_waddr, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_executeUnit_flush, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_executeUnit_allow_to_go, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_executeUnit_do_flush, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_executeUnit_fu_allow_to_go, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_executeUnit_fu_stall, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_memoryUnit_flush, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_memoryUnit_mem_stall, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_memoryUnit_allow_to_go, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_memoryUnit_do_flush, // @[playground/src/ctrl/Ctrl.scala 10:14]
  input        io_memoryUnit_complete_single_request, // @[playground/src/ctrl/Ctrl.scala 10:14]
  output       io_writeBackUnit_allow_to_go // @[playground/src/ctrl/Ctrl.scala 10:14]
);
  wire  _inst0_lw_stall_T_5 = io_decodeUnit_inst0_src2_ren & io_decodeUnit_inst0_src2_raddr ==
    io_executeUnit_inst_0_reg_waddr; // @[playground/src/ctrl/Ctrl.scala 21:36]
  wire  _inst0_lw_stall_T_6 = io_decodeUnit_inst0_src1_ren & io_decodeUnit_inst0_src1_raddr ==
    io_executeUnit_inst_0_reg_waddr | _inst0_lw_stall_T_5; // @[playground/src/ctrl/Ctrl.scala 20:106]
  wire  inst0_lw_stall = io_executeUnit_inst_0_is_load & |io_executeUnit_inst_0_reg_waddr & _inst0_lw_stall_T_6; // @[playground/src/ctrl/Ctrl.scala 19:97]
  wire  _inst1_lw_stall_T_5 = io_decodeUnit_inst0_src2_ren & io_decodeUnit_inst0_src2_raddr ==
    io_executeUnit_inst_1_reg_waddr; // @[playground/src/ctrl/Ctrl.scala 24:36]
  wire  _inst1_lw_stall_T_6 = io_decodeUnit_inst0_src1_ren & io_decodeUnit_inst0_src1_raddr ==
    io_executeUnit_inst_1_reg_waddr | _inst1_lw_stall_T_5; // @[playground/src/ctrl/Ctrl.scala 23:106]
  wire  inst1_lw_stall = io_executeUnit_inst_1_is_load & |io_executeUnit_inst_1_reg_waddr & _inst1_lw_stall_T_6; // @[playground/src/ctrl/Ctrl.scala 22:97]
  wire  lw_stall = inst0_lw_stall | inst1_lw_stall; // @[playground/src/ctrl/Ctrl.scala 25:33]
  wire  longest_stall = io_executeUnit_fu_stall | io_cacheCtrl_iCache_stall | io_memoryUnit_mem_stall; // @[playground/src/ctrl/Ctrl.scala 27:58]
  assign io_fetchUnit_allow_to_go = ~io_cacheCtrl_iCache_stall; // @[playground/src/ctrl/Ctrl.scala 29:35]
  assign io_decodeUnit_allow_to_go = ~(lw_stall | longest_stall); // @[playground/src/ctrl/Ctrl.scala 30:35]
  assign io_decodeUnit_do_flush = io_memoryUnit_flush | io_executeUnit_flush | io_decodeUnit_branch; // @[playground/src/ctrl/Ctrl.scala 36:76]
  assign io_executeUnit_allow_to_go = ~longest_stall; // @[playground/src/ctrl/Ctrl.scala 31:35]
  assign io_executeUnit_do_flush = io_memoryUnit_flush | io_executeUnit_flush; // @[playground/src/ctrl/Ctrl.scala 37:52]
  assign io_executeUnit_fu_allow_to_go = io_memoryUnit_allow_to_go; // @[playground/src/ctrl/Ctrl.scala 41:33]
  assign io_memoryUnit_allow_to_go = ~longest_stall; // @[playground/src/ctrl/Ctrl.scala 32:35]
  assign io_memoryUnit_do_flush = io_memoryUnit_flush; // @[playground/src/ctrl/Ctrl.scala 38:29]
  assign io_writeBackUnit_allow_to_go = ~longest_stall; // @[playground/src/ctrl/Ctrl.scala 33:35]
endmodule
module FetchUnit(
  input         clock,
  input         reset,
  input         io_memory_flush, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input  [63:0] io_memory_target, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input         io_decode_branch, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input  [63:0] io_decode_target, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input         io_execute_flush, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input  [63:0] io_execute_target, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input         io_instFifo_full, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input         io_iCache_inst_valid_0, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  input         io_iCache_inst_valid_1, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  output [63:0] io_iCache_pc, // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
  output [63:0] io_iCache_pc_next // @[playground/src/pipeline/fetch/FetchUnit.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] pc; // @[playground/src/pipeline/fetch/FetchUnit.scala 35:19]
  wire [63:0] _pc_next_temp_T_1 = pc + 64'h4; // @[playground/src/pipeline/fetch/FetchUnit.scala 45:26]
  wire [63:0] _GEN_0 = io_iCache_inst_valid_0 ? _pc_next_temp_T_1 : pc; // @[playground/src/pipeline/fetch/FetchUnit.scala 42:16 44:35 45:20]
  wire [63:0] _pc_next_temp_T_3 = pc + 64'h8; // @[playground/src/pipeline/fetch/FetchUnit.scala 45:26]
  wire [63:0] pc_next_temp = io_iCache_inst_valid_1 ? _pc_next_temp_T_3 : _GEN_0; // @[playground/src/pipeline/fetch/FetchUnit.scala 44:35 45:20]
  wire [63:0] _io_iCache_pc_next_T = io_instFifo_full ? pc : pc_next_temp; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _io_iCache_pc_next_T_1 = io_decode_branch ? io_decode_target : _io_iCache_pc_next_T; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _io_iCache_pc_next_T_2 = io_execute_flush ? io_execute_target : _io_iCache_pc_next_T_1; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_iCache_pc = pc; // @[playground/src/pipeline/fetch/FetchUnit.scala 36:16]
  assign io_iCache_pc_next = io_memory_flush ? io_memory_target : _io_iCache_pc_next_T_2; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/fetch/FetchUnit.scala 35:19]
      pc <= 64'h80000000; // @[playground/src/pipeline/fetch/FetchUnit.scala 35:19]
    end else begin
      pc <= io_iCache_pc_next; // @[playground/src/pipeline/fetch/FetchUnit.scala 35:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AdaptiveTwoLevelPredictor(
  input         clock,
  input         reset,
  input  [63:0] io_decode_pc, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input         io_decode_info_valid, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [2:0]  io_decode_info_fusel, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [6:0]  io_decode_info_op, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [63:0] io_decode_info_imm, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [5:0]  io_decode_pht_index, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  output        io_decode_branch_inst, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  output        io_decode_branch, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  output [63:0] io_decode_target, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  output [5:0]  io_decode_update_pht_index, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [63:0] io_instBuffer_pc_0, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [63:0] io_instBuffer_pc_1, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  output [5:0]  io_instBuffer_pht_index_0, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  output [5:0]  io_instBuffer_pht_index_1, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [63:0] io_execute_pc, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input  [5:0]  io_execute_update_pht_index, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input         io_execute_branch_inst, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
  input         io_execute_branch // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 107:21]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
`endif // RANDOMIZE_REG_INIT
  wire  _io_decode_branch_inst_T = 3'h5 == io_decode_info_fusel; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 114:16]
  wire  _io_decode_branch_inst_T_1 = io_decode_info_valid & _io_decode_branch_inst_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 113:49]
  wire  _io_decode_branch_inst_T_3 = ~io_decode_info_op[3]; // @[playground/src/defines/isa/Instructions.scala 74:36]
  reg [5:0] bht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [5:0] bht_31; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
  reg [1:0] pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_31; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_32; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_33; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_34; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_35; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_36; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_37; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_38; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_39; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_40; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_41; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_42; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_43; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_44; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_45; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_46; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_47; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_48; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_49; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_50; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_51; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_52; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_53; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_54; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_55; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_56; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_57; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_58; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_59; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_60; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_61; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_62; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  reg [1:0] pht_63; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
  wire [5:0] _GEN_1 = 5'h1 == io_instBuffer_pc_0[6:2] ? bht_1 : bht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_2 = 5'h2 == io_instBuffer_pc_0[6:2] ? bht_2 : _GEN_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_3 = 5'h3 == io_instBuffer_pc_0[6:2] ? bht_3 : _GEN_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_4 = 5'h4 == io_instBuffer_pc_0[6:2] ? bht_4 : _GEN_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_5 = 5'h5 == io_instBuffer_pc_0[6:2] ? bht_5 : _GEN_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_6 = 5'h6 == io_instBuffer_pc_0[6:2] ? bht_6 : _GEN_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_7 = 5'h7 == io_instBuffer_pc_0[6:2] ? bht_7 : _GEN_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_8 = 5'h8 == io_instBuffer_pc_0[6:2] ? bht_8 : _GEN_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_9 = 5'h9 == io_instBuffer_pc_0[6:2] ? bht_9 : _GEN_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_10 = 5'ha == io_instBuffer_pc_0[6:2] ? bht_10 : _GEN_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_11 = 5'hb == io_instBuffer_pc_0[6:2] ? bht_11 : _GEN_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_12 = 5'hc == io_instBuffer_pc_0[6:2] ? bht_12 : _GEN_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_13 = 5'hd == io_instBuffer_pc_0[6:2] ? bht_13 : _GEN_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_14 = 5'he == io_instBuffer_pc_0[6:2] ? bht_14 : _GEN_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_15 = 5'hf == io_instBuffer_pc_0[6:2] ? bht_15 : _GEN_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_16 = 5'h10 == io_instBuffer_pc_0[6:2] ? bht_16 : _GEN_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_17 = 5'h11 == io_instBuffer_pc_0[6:2] ? bht_17 : _GEN_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_18 = 5'h12 == io_instBuffer_pc_0[6:2] ? bht_18 : _GEN_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_19 = 5'h13 == io_instBuffer_pc_0[6:2] ? bht_19 : _GEN_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_20 = 5'h14 == io_instBuffer_pc_0[6:2] ? bht_20 : _GEN_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_21 = 5'h15 == io_instBuffer_pc_0[6:2] ? bht_21 : _GEN_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_22 = 5'h16 == io_instBuffer_pc_0[6:2] ? bht_22 : _GEN_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_23 = 5'h17 == io_instBuffer_pc_0[6:2] ? bht_23 : _GEN_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_24 = 5'h18 == io_instBuffer_pc_0[6:2] ? bht_24 : _GEN_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_25 = 5'h19 == io_instBuffer_pc_0[6:2] ? bht_25 : _GEN_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_26 = 5'h1a == io_instBuffer_pc_0[6:2] ? bht_26 : _GEN_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_27 = 5'h1b == io_instBuffer_pc_0[6:2] ? bht_27 : _GEN_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_28 = 5'h1c == io_instBuffer_pc_0[6:2] ? bht_28 : _GEN_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_29 = 5'h1d == io_instBuffer_pc_0[6:2] ? bht_29 : _GEN_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_30 = 5'h1e == io_instBuffer_pc_0[6:2] ? bht_30 : _GEN_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_33 = 5'h1 == io_instBuffer_pc_1[6:2] ? bht_1 : bht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_34 = 5'h2 == io_instBuffer_pc_1[6:2] ? bht_2 : _GEN_33; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_35 = 5'h3 == io_instBuffer_pc_1[6:2] ? bht_3 : _GEN_34; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_36 = 5'h4 == io_instBuffer_pc_1[6:2] ? bht_4 : _GEN_35; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_37 = 5'h5 == io_instBuffer_pc_1[6:2] ? bht_5 : _GEN_36; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_38 = 5'h6 == io_instBuffer_pc_1[6:2] ? bht_6 : _GEN_37; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_39 = 5'h7 == io_instBuffer_pc_1[6:2] ? bht_7 : _GEN_38; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_40 = 5'h8 == io_instBuffer_pc_1[6:2] ? bht_8 : _GEN_39; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_41 = 5'h9 == io_instBuffer_pc_1[6:2] ? bht_9 : _GEN_40; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_42 = 5'ha == io_instBuffer_pc_1[6:2] ? bht_10 : _GEN_41; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_43 = 5'hb == io_instBuffer_pc_1[6:2] ? bht_11 : _GEN_42; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_44 = 5'hc == io_instBuffer_pc_1[6:2] ? bht_12 : _GEN_43; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_45 = 5'hd == io_instBuffer_pc_1[6:2] ? bht_13 : _GEN_44; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_46 = 5'he == io_instBuffer_pc_1[6:2] ? bht_14 : _GEN_45; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_47 = 5'hf == io_instBuffer_pc_1[6:2] ? bht_15 : _GEN_46; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_48 = 5'h10 == io_instBuffer_pc_1[6:2] ? bht_16 : _GEN_47; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_49 = 5'h11 == io_instBuffer_pc_1[6:2] ? bht_17 : _GEN_48; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_50 = 5'h12 == io_instBuffer_pc_1[6:2] ? bht_18 : _GEN_49; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_51 = 5'h13 == io_instBuffer_pc_1[6:2] ? bht_19 : _GEN_50; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_52 = 5'h14 == io_instBuffer_pc_1[6:2] ? bht_20 : _GEN_51; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_53 = 5'h15 == io_instBuffer_pc_1[6:2] ? bht_21 : _GEN_52; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_54 = 5'h16 == io_instBuffer_pc_1[6:2] ? bht_22 : _GEN_53; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_55 = 5'h17 == io_instBuffer_pc_1[6:2] ? bht_23 : _GEN_54; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_56 = 5'h18 == io_instBuffer_pc_1[6:2] ? bht_24 : _GEN_55; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_57 = 5'h19 == io_instBuffer_pc_1[6:2] ? bht_25 : _GEN_56; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_58 = 5'h1a == io_instBuffer_pc_1[6:2] ? bht_26 : _GEN_57; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_59 = 5'h1b == io_instBuffer_pc_1[6:2] ? bht_27 : _GEN_58; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_60 = 5'h1c == io_instBuffer_pc_1[6:2] ? bht_28 : _GEN_59; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_61 = 5'h1d == io_instBuffer_pc_1[6:2] ? bht_29 : _GEN_60; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [5:0] _GEN_62 = 5'h1e == io_instBuffer_pc_1[6:2] ? bht_30 : _GEN_61; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  wire [1:0] _GEN_65 = 6'h1 == io_decode_pht_index ? pht_1 : pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_66 = 6'h2 == io_decode_pht_index ? pht_2 : _GEN_65; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_67 = 6'h3 == io_decode_pht_index ? pht_3 : _GEN_66; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_68 = 6'h4 == io_decode_pht_index ? pht_4 : _GEN_67; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_69 = 6'h5 == io_decode_pht_index ? pht_5 : _GEN_68; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_70 = 6'h6 == io_decode_pht_index ? pht_6 : _GEN_69; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_71 = 6'h7 == io_decode_pht_index ? pht_7 : _GEN_70; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_72 = 6'h8 == io_decode_pht_index ? pht_8 : _GEN_71; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_73 = 6'h9 == io_decode_pht_index ? pht_9 : _GEN_72; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_74 = 6'ha == io_decode_pht_index ? pht_10 : _GEN_73; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_75 = 6'hb == io_decode_pht_index ? pht_11 : _GEN_74; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_76 = 6'hc == io_decode_pht_index ? pht_12 : _GEN_75; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_77 = 6'hd == io_decode_pht_index ? pht_13 : _GEN_76; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_78 = 6'he == io_decode_pht_index ? pht_14 : _GEN_77; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_79 = 6'hf == io_decode_pht_index ? pht_15 : _GEN_78; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_80 = 6'h10 == io_decode_pht_index ? pht_16 : _GEN_79; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_81 = 6'h11 == io_decode_pht_index ? pht_17 : _GEN_80; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_82 = 6'h12 == io_decode_pht_index ? pht_18 : _GEN_81; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_83 = 6'h13 == io_decode_pht_index ? pht_19 : _GEN_82; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_84 = 6'h14 == io_decode_pht_index ? pht_20 : _GEN_83; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_85 = 6'h15 == io_decode_pht_index ? pht_21 : _GEN_84; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_86 = 6'h16 == io_decode_pht_index ? pht_22 : _GEN_85; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_87 = 6'h17 == io_decode_pht_index ? pht_23 : _GEN_86; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_88 = 6'h18 == io_decode_pht_index ? pht_24 : _GEN_87; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_89 = 6'h19 == io_decode_pht_index ? pht_25 : _GEN_88; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_90 = 6'h1a == io_decode_pht_index ? pht_26 : _GEN_89; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_91 = 6'h1b == io_decode_pht_index ? pht_27 : _GEN_90; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_92 = 6'h1c == io_decode_pht_index ? pht_28 : _GEN_91; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_93 = 6'h1d == io_decode_pht_index ? pht_29 : _GEN_92; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_94 = 6'h1e == io_decode_pht_index ? pht_30 : _GEN_93; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_95 = 6'h1f == io_decode_pht_index ? pht_31 : _GEN_94; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_96 = 6'h20 == io_decode_pht_index ? pht_32 : _GEN_95; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_97 = 6'h21 == io_decode_pht_index ? pht_33 : _GEN_96; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_98 = 6'h22 == io_decode_pht_index ? pht_34 : _GEN_97; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_99 = 6'h23 == io_decode_pht_index ? pht_35 : _GEN_98; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_100 = 6'h24 == io_decode_pht_index ? pht_36 : _GEN_99; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_101 = 6'h25 == io_decode_pht_index ? pht_37 : _GEN_100; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_102 = 6'h26 == io_decode_pht_index ? pht_38 : _GEN_101; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_103 = 6'h27 == io_decode_pht_index ? pht_39 : _GEN_102; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_104 = 6'h28 == io_decode_pht_index ? pht_40 : _GEN_103; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_105 = 6'h29 == io_decode_pht_index ? pht_41 : _GEN_104; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_106 = 6'h2a == io_decode_pht_index ? pht_42 : _GEN_105; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_107 = 6'h2b == io_decode_pht_index ? pht_43 : _GEN_106; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_108 = 6'h2c == io_decode_pht_index ? pht_44 : _GEN_107; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_109 = 6'h2d == io_decode_pht_index ? pht_45 : _GEN_108; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_110 = 6'h2e == io_decode_pht_index ? pht_46 : _GEN_109; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_111 = 6'h2f == io_decode_pht_index ? pht_47 : _GEN_110; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_112 = 6'h30 == io_decode_pht_index ? pht_48 : _GEN_111; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_113 = 6'h31 == io_decode_pht_index ? pht_49 : _GEN_112; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_114 = 6'h32 == io_decode_pht_index ? pht_50 : _GEN_113; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_115 = 6'h33 == io_decode_pht_index ? pht_51 : _GEN_114; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_116 = 6'h34 == io_decode_pht_index ? pht_52 : _GEN_115; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_117 = 6'h35 == io_decode_pht_index ? pht_53 : _GEN_116; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_118 = 6'h36 == io_decode_pht_index ? pht_54 : _GEN_117; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_119 = 6'h37 == io_decode_pht_index ? pht_55 : _GEN_118; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_120 = 6'h38 == io_decode_pht_index ? pht_56 : _GEN_119; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_121 = 6'h39 == io_decode_pht_index ? pht_57 : _GEN_120; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_122 = 6'h3a == io_decode_pht_index ? pht_58 : _GEN_121; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_123 = 6'h3b == io_decode_pht_index ? pht_59 : _GEN_122; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_124 = 6'h3c == io_decode_pht_index ? pht_60 : _GEN_123; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_125 = 6'h3d == io_decode_pht_index ? pht_61 : _GEN_124; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_126 = 6'h3e == io_decode_pht_index ? pht_62 : _GEN_125; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [1:0] _GEN_127 = 6'h3f == io_decode_pht_index ? pht_63 : _GEN_126; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:{46,46}]
  wire [5:0] _GEN_129 = 5'h1 == io_decode_pc[6:2] ? bht_1 : bht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_130 = 5'h2 == io_decode_pc[6:2] ? bht_2 : _GEN_129; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_131 = 5'h3 == io_decode_pc[6:2] ? bht_3 : _GEN_130; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_132 = 5'h4 == io_decode_pc[6:2] ? bht_4 : _GEN_131; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_133 = 5'h5 == io_decode_pc[6:2] ? bht_5 : _GEN_132; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_134 = 5'h6 == io_decode_pc[6:2] ? bht_6 : _GEN_133; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_135 = 5'h7 == io_decode_pc[6:2] ? bht_7 : _GEN_134; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_136 = 5'h8 == io_decode_pc[6:2] ? bht_8 : _GEN_135; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_137 = 5'h9 == io_decode_pc[6:2] ? bht_9 : _GEN_136; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_138 = 5'ha == io_decode_pc[6:2] ? bht_10 : _GEN_137; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_139 = 5'hb == io_decode_pc[6:2] ? bht_11 : _GEN_138; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_140 = 5'hc == io_decode_pc[6:2] ? bht_12 : _GEN_139; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_141 = 5'hd == io_decode_pc[6:2] ? bht_13 : _GEN_140; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_142 = 5'he == io_decode_pc[6:2] ? bht_14 : _GEN_141; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_143 = 5'hf == io_decode_pc[6:2] ? bht_15 : _GEN_142; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_144 = 5'h10 == io_decode_pc[6:2] ? bht_16 : _GEN_143; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_145 = 5'h11 == io_decode_pc[6:2] ? bht_17 : _GEN_144; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_146 = 5'h12 == io_decode_pc[6:2] ? bht_18 : _GEN_145; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_147 = 5'h13 == io_decode_pc[6:2] ? bht_19 : _GEN_146; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_148 = 5'h14 == io_decode_pc[6:2] ? bht_20 : _GEN_147; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_149 = 5'h15 == io_decode_pc[6:2] ? bht_21 : _GEN_148; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_150 = 5'h16 == io_decode_pc[6:2] ? bht_22 : _GEN_149; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_151 = 5'h17 == io_decode_pc[6:2] ? bht_23 : _GEN_150; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_152 = 5'h18 == io_decode_pc[6:2] ? bht_24 : _GEN_151; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_153 = 5'h19 == io_decode_pc[6:2] ? bht_25 : _GEN_152; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_154 = 5'h1a == io_decode_pc[6:2] ? bht_26 : _GEN_153; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_155 = 5'h1b == io_decode_pc[6:2] ? bht_27 : _GEN_154; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_156 = 5'h1c == io_decode_pc[6:2] ? bht_28 : _GEN_155; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_157 = 5'h1d == io_decode_pc[6:2] ? bht_29 : _GEN_156; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [5:0] _GEN_158 = 5'h1e == io_decode_pc[6:2] ? bht_30 : _GEN_157; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  wire [4:0] update_bht_index = io_execute_pc[6:2]; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 129:39]
  wire [5:0] _GEN_161 = 5'h1 == update_bht_index ? bht_1 : bht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_162 = 5'h2 == update_bht_index ? bht_2 : _GEN_161; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_163 = 5'h3 == update_bht_index ? bht_3 : _GEN_162; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_164 = 5'h4 == update_bht_index ? bht_4 : _GEN_163; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_165 = 5'h5 == update_bht_index ? bht_5 : _GEN_164; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_166 = 5'h6 == update_bht_index ? bht_6 : _GEN_165; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_167 = 5'h7 == update_bht_index ? bht_7 : _GEN_166; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_168 = 5'h8 == update_bht_index ? bht_8 : _GEN_167; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_169 = 5'h9 == update_bht_index ? bht_9 : _GEN_168; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_170 = 5'ha == update_bht_index ? bht_10 : _GEN_169; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_171 = 5'hb == update_bht_index ? bht_11 : _GEN_170; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_172 = 5'hc == update_bht_index ? bht_12 : _GEN_171; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_173 = 5'hd == update_bht_index ? bht_13 : _GEN_172; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_174 = 5'he == update_bht_index ? bht_14 : _GEN_173; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_175 = 5'hf == update_bht_index ? bht_15 : _GEN_174; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_176 = 5'h10 == update_bht_index ? bht_16 : _GEN_175; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_177 = 5'h11 == update_bht_index ? bht_17 : _GEN_176; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_178 = 5'h12 == update_bht_index ? bht_18 : _GEN_177; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_179 = 5'h13 == update_bht_index ? bht_19 : _GEN_178; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_180 = 5'h14 == update_bht_index ? bht_20 : _GEN_179; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_181 = 5'h15 == update_bht_index ? bht_21 : _GEN_180; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_182 = 5'h16 == update_bht_index ? bht_22 : _GEN_181; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_183 = 5'h17 == update_bht_index ? bht_23 : _GEN_182; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_184 = 5'h18 == update_bht_index ? bht_24 : _GEN_183; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_185 = 5'h19 == update_bht_index ? bht_25 : _GEN_184; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_186 = 5'h1a == update_bht_index ? bht_26 : _GEN_185; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_187 = 5'h1b == update_bht_index ? bht_27 : _GEN_186; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_188 = 5'h1c == update_bht_index ? bht_28 : _GEN_187; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_189 = 5'h1d == update_bht_index ? bht_29 : _GEN_188; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_190 = 5'h1e == update_bht_index ? bht_30 : _GEN_189; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _GEN_191 = 5'h1f == update_bht_index ? bht_31 : _GEN_190; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:{55,55}]
  wire [5:0] _bht_T_1 = {_GEN_191[4:0],io_execute_branch}; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:33]
  wire [1:0] _GEN_225 = 6'h1 == io_execute_update_pht_index ? pht_1 : pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_226 = 6'h2 == io_execute_update_pht_index ? pht_2 : _GEN_225; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_227 = 6'h3 == io_execute_update_pht_index ? pht_3 : _GEN_226; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_228 = 6'h4 == io_execute_update_pht_index ? pht_4 : _GEN_227; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_229 = 6'h5 == io_execute_update_pht_index ? pht_5 : _GEN_228; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_230 = 6'h6 == io_execute_update_pht_index ? pht_6 : _GEN_229; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_231 = 6'h7 == io_execute_update_pht_index ? pht_7 : _GEN_230; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_232 = 6'h8 == io_execute_update_pht_index ? pht_8 : _GEN_231; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_233 = 6'h9 == io_execute_update_pht_index ? pht_9 : _GEN_232; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_234 = 6'ha == io_execute_update_pht_index ? pht_10 : _GEN_233; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_235 = 6'hb == io_execute_update_pht_index ? pht_11 : _GEN_234; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_236 = 6'hc == io_execute_update_pht_index ? pht_12 : _GEN_235; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_237 = 6'hd == io_execute_update_pht_index ? pht_13 : _GEN_236; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_238 = 6'he == io_execute_update_pht_index ? pht_14 : _GEN_237; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_239 = 6'hf == io_execute_update_pht_index ? pht_15 : _GEN_238; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_240 = 6'h10 == io_execute_update_pht_index ? pht_16 : _GEN_239; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_241 = 6'h11 == io_execute_update_pht_index ? pht_17 : _GEN_240; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_242 = 6'h12 == io_execute_update_pht_index ? pht_18 : _GEN_241; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_243 = 6'h13 == io_execute_update_pht_index ? pht_19 : _GEN_242; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_244 = 6'h14 == io_execute_update_pht_index ? pht_20 : _GEN_243; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_245 = 6'h15 == io_execute_update_pht_index ? pht_21 : _GEN_244; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_246 = 6'h16 == io_execute_update_pht_index ? pht_22 : _GEN_245; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_247 = 6'h17 == io_execute_update_pht_index ? pht_23 : _GEN_246; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_248 = 6'h18 == io_execute_update_pht_index ? pht_24 : _GEN_247; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_249 = 6'h19 == io_execute_update_pht_index ? pht_25 : _GEN_248; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_250 = 6'h1a == io_execute_update_pht_index ? pht_26 : _GEN_249; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_251 = 6'h1b == io_execute_update_pht_index ? pht_27 : _GEN_250; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_252 = 6'h1c == io_execute_update_pht_index ? pht_28 : _GEN_251; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_253 = 6'h1d == io_execute_update_pht_index ? pht_29 : _GEN_252; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_254 = 6'h1e == io_execute_update_pht_index ? pht_30 : _GEN_253; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_255 = 6'h1f == io_execute_update_pht_index ? pht_31 : _GEN_254; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_256 = 6'h20 == io_execute_update_pht_index ? pht_32 : _GEN_255; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_257 = 6'h21 == io_execute_update_pht_index ? pht_33 : _GEN_256; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_258 = 6'h22 == io_execute_update_pht_index ? pht_34 : _GEN_257; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_259 = 6'h23 == io_execute_update_pht_index ? pht_35 : _GEN_258; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_260 = 6'h24 == io_execute_update_pht_index ? pht_36 : _GEN_259; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_261 = 6'h25 == io_execute_update_pht_index ? pht_37 : _GEN_260; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_262 = 6'h26 == io_execute_update_pht_index ? pht_38 : _GEN_261; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_263 = 6'h27 == io_execute_update_pht_index ? pht_39 : _GEN_262; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_264 = 6'h28 == io_execute_update_pht_index ? pht_40 : _GEN_263; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_265 = 6'h29 == io_execute_update_pht_index ? pht_41 : _GEN_264; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_266 = 6'h2a == io_execute_update_pht_index ? pht_42 : _GEN_265; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_267 = 6'h2b == io_execute_update_pht_index ? pht_43 : _GEN_266; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_268 = 6'h2c == io_execute_update_pht_index ? pht_44 : _GEN_267; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_269 = 6'h2d == io_execute_update_pht_index ? pht_45 : _GEN_268; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_270 = 6'h2e == io_execute_update_pht_index ? pht_46 : _GEN_269; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_271 = 6'h2f == io_execute_update_pht_index ? pht_47 : _GEN_270; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_272 = 6'h30 == io_execute_update_pht_index ? pht_48 : _GEN_271; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_273 = 6'h31 == io_execute_update_pht_index ? pht_49 : _GEN_272; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_274 = 6'h32 == io_execute_update_pht_index ? pht_50 : _GEN_273; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_275 = 6'h33 == io_execute_update_pht_index ? pht_51 : _GEN_274; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_276 = 6'h34 == io_execute_update_pht_index ? pht_52 : _GEN_275; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_277 = 6'h35 == io_execute_update_pht_index ? pht_53 : _GEN_276; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_278 = 6'h36 == io_execute_update_pht_index ? pht_54 : _GEN_277; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_279 = 6'h37 == io_execute_update_pht_index ? pht_55 : _GEN_278; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_280 = 6'h38 == io_execute_update_pht_index ? pht_56 : _GEN_279; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_281 = 6'h39 == io_execute_update_pht_index ? pht_57 : _GEN_280; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_282 = 6'h3a == io_execute_update_pht_index ? pht_58 : _GEN_281; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_283 = 6'h3b == io_execute_update_pht_index ? pht_59 : _GEN_282; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_284 = 6'h3c == io_execute_update_pht_index ? pht_60 : _GEN_283; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_285 = 6'h3d == io_execute_update_pht_index ? pht_61 : _GEN_284; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_286 = 6'h3e == io_execute_update_pht_index ? pht_62 : _GEN_285; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _GEN_287 = 6'h3f == io_execute_update_pht_index ? pht_63 : _GEN_286; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:{35,35}]
  wire [1:0] _pht_T = io_execute_branch ? 2'h1 : 2'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:37]
  wire [1:0] _pht_T_1 = io_execute_branch ? 2'h2 : 2'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 139:37]
  wire [1:0] _GEN_352 = 6'h0 == io_execute_update_pht_index ? _pht_T_1 : pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_353 = 6'h1 == io_execute_update_pht_index ? _pht_T_1 : pht_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_354 = 6'h2 == io_execute_update_pht_index ? _pht_T_1 : pht_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_355 = 6'h3 == io_execute_update_pht_index ? _pht_T_1 : pht_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_356 = 6'h4 == io_execute_update_pht_index ? _pht_T_1 : pht_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_357 = 6'h5 == io_execute_update_pht_index ? _pht_T_1 : pht_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_358 = 6'h6 == io_execute_update_pht_index ? _pht_T_1 : pht_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_359 = 6'h7 == io_execute_update_pht_index ? _pht_T_1 : pht_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_360 = 6'h8 == io_execute_update_pht_index ? _pht_T_1 : pht_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_361 = 6'h9 == io_execute_update_pht_index ? _pht_T_1 : pht_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_362 = 6'ha == io_execute_update_pht_index ? _pht_T_1 : pht_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_363 = 6'hb == io_execute_update_pht_index ? _pht_T_1 : pht_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_364 = 6'hc == io_execute_update_pht_index ? _pht_T_1 : pht_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_365 = 6'hd == io_execute_update_pht_index ? _pht_T_1 : pht_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_366 = 6'he == io_execute_update_pht_index ? _pht_T_1 : pht_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_367 = 6'hf == io_execute_update_pht_index ? _pht_T_1 : pht_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_368 = 6'h10 == io_execute_update_pht_index ? _pht_T_1 : pht_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_369 = 6'h11 == io_execute_update_pht_index ? _pht_T_1 : pht_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_370 = 6'h12 == io_execute_update_pht_index ? _pht_T_1 : pht_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_371 = 6'h13 == io_execute_update_pht_index ? _pht_T_1 : pht_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_372 = 6'h14 == io_execute_update_pht_index ? _pht_T_1 : pht_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_373 = 6'h15 == io_execute_update_pht_index ? _pht_T_1 : pht_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_374 = 6'h16 == io_execute_update_pht_index ? _pht_T_1 : pht_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_375 = 6'h17 == io_execute_update_pht_index ? _pht_T_1 : pht_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_376 = 6'h18 == io_execute_update_pht_index ? _pht_T_1 : pht_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_377 = 6'h19 == io_execute_update_pht_index ? _pht_T_1 : pht_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_378 = 6'h1a == io_execute_update_pht_index ? _pht_T_1 : pht_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_379 = 6'h1b == io_execute_update_pht_index ? _pht_T_1 : pht_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_380 = 6'h1c == io_execute_update_pht_index ? _pht_T_1 : pht_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_381 = 6'h1d == io_execute_update_pht_index ? _pht_T_1 : pht_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_382 = 6'h1e == io_execute_update_pht_index ? _pht_T_1 : pht_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_383 = 6'h1f == io_execute_update_pht_index ? _pht_T_1 : pht_31; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_384 = 6'h20 == io_execute_update_pht_index ? _pht_T_1 : pht_32; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_385 = 6'h21 == io_execute_update_pht_index ? _pht_T_1 : pht_33; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_386 = 6'h22 == io_execute_update_pht_index ? _pht_T_1 : pht_34; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_387 = 6'h23 == io_execute_update_pht_index ? _pht_T_1 : pht_35; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_388 = 6'h24 == io_execute_update_pht_index ? _pht_T_1 : pht_36; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_389 = 6'h25 == io_execute_update_pht_index ? _pht_T_1 : pht_37; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_390 = 6'h26 == io_execute_update_pht_index ? _pht_T_1 : pht_38; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_391 = 6'h27 == io_execute_update_pht_index ? _pht_T_1 : pht_39; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_392 = 6'h28 == io_execute_update_pht_index ? _pht_T_1 : pht_40; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_393 = 6'h29 == io_execute_update_pht_index ? _pht_T_1 : pht_41; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_394 = 6'h2a == io_execute_update_pht_index ? _pht_T_1 : pht_42; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_395 = 6'h2b == io_execute_update_pht_index ? _pht_T_1 : pht_43; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_396 = 6'h2c == io_execute_update_pht_index ? _pht_T_1 : pht_44; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_397 = 6'h2d == io_execute_update_pht_index ? _pht_T_1 : pht_45; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_398 = 6'h2e == io_execute_update_pht_index ? _pht_T_1 : pht_46; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_399 = 6'h2f == io_execute_update_pht_index ? _pht_T_1 : pht_47; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_400 = 6'h30 == io_execute_update_pht_index ? _pht_T_1 : pht_48; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_401 = 6'h31 == io_execute_update_pht_index ? _pht_T_1 : pht_49; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_402 = 6'h32 == io_execute_update_pht_index ? _pht_T_1 : pht_50; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_403 = 6'h33 == io_execute_update_pht_index ? _pht_T_1 : pht_51; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_404 = 6'h34 == io_execute_update_pht_index ? _pht_T_1 : pht_52; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_405 = 6'h35 == io_execute_update_pht_index ? _pht_T_1 : pht_53; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_406 = 6'h36 == io_execute_update_pht_index ? _pht_T_1 : pht_54; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_407 = 6'h37 == io_execute_update_pht_index ? _pht_T_1 : pht_55; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_408 = 6'h38 == io_execute_update_pht_index ? _pht_T_1 : pht_56; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_409 = 6'h39 == io_execute_update_pht_index ? _pht_T_1 : pht_57; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_410 = 6'h3a == io_execute_update_pht_index ? _pht_T_1 : pht_58; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_411 = 6'h3b == io_execute_update_pht_index ? _pht_T_1 : pht_59; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_412 = 6'h3c == io_execute_update_pht_index ? _pht_T_1 : pht_60; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_413 = 6'h3d == io_execute_update_pht_index ? _pht_T_1 : pht_61; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_414 = 6'h3e == io_execute_update_pht_index ? _pht_T_1 : pht_62; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _GEN_415 = 6'h3f == io_execute_update_pht_index ? _pht_T_1 : pht_63; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 139:{31,31}]
  wire [1:0] _pht_T_2 = io_execute_branch ? 2'h3 : 2'h1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 142:37]
  wire [1:0] _GEN_416 = 6'h0 == io_execute_update_pht_index ? _pht_T_2 : pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_417 = 6'h1 == io_execute_update_pht_index ? _pht_T_2 : pht_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_418 = 6'h2 == io_execute_update_pht_index ? _pht_T_2 : pht_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_419 = 6'h3 == io_execute_update_pht_index ? _pht_T_2 : pht_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_420 = 6'h4 == io_execute_update_pht_index ? _pht_T_2 : pht_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_421 = 6'h5 == io_execute_update_pht_index ? _pht_T_2 : pht_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_422 = 6'h6 == io_execute_update_pht_index ? _pht_T_2 : pht_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_423 = 6'h7 == io_execute_update_pht_index ? _pht_T_2 : pht_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_424 = 6'h8 == io_execute_update_pht_index ? _pht_T_2 : pht_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_425 = 6'h9 == io_execute_update_pht_index ? _pht_T_2 : pht_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_426 = 6'ha == io_execute_update_pht_index ? _pht_T_2 : pht_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_427 = 6'hb == io_execute_update_pht_index ? _pht_T_2 : pht_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_428 = 6'hc == io_execute_update_pht_index ? _pht_T_2 : pht_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_429 = 6'hd == io_execute_update_pht_index ? _pht_T_2 : pht_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_430 = 6'he == io_execute_update_pht_index ? _pht_T_2 : pht_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_431 = 6'hf == io_execute_update_pht_index ? _pht_T_2 : pht_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_432 = 6'h10 == io_execute_update_pht_index ? _pht_T_2 : pht_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_433 = 6'h11 == io_execute_update_pht_index ? _pht_T_2 : pht_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_434 = 6'h12 == io_execute_update_pht_index ? _pht_T_2 : pht_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_435 = 6'h13 == io_execute_update_pht_index ? _pht_T_2 : pht_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_436 = 6'h14 == io_execute_update_pht_index ? _pht_T_2 : pht_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_437 = 6'h15 == io_execute_update_pht_index ? _pht_T_2 : pht_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_438 = 6'h16 == io_execute_update_pht_index ? _pht_T_2 : pht_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_439 = 6'h17 == io_execute_update_pht_index ? _pht_T_2 : pht_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_440 = 6'h18 == io_execute_update_pht_index ? _pht_T_2 : pht_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_441 = 6'h19 == io_execute_update_pht_index ? _pht_T_2 : pht_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_442 = 6'h1a == io_execute_update_pht_index ? _pht_T_2 : pht_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_443 = 6'h1b == io_execute_update_pht_index ? _pht_T_2 : pht_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_444 = 6'h1c == io_execute_update_pht_index ? _pht_T_2 : pht_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_445 = 6'h1d == io_execute_update_pht_index ? _pht_T_2 : pht_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_446 = 6'h1e == io_execute_update_pht_index ? _pht_T_2 : pht_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_447 = 6'h1f == io_execute_update_pht_index ? _pht_T_2 : pht_31; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_448 = 6'h20 == io_execute_update_pht_index ? _pht_T_2 : pht_32; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_449 = 6'h21 == io_execute_update_pht_index ? _pht_T_2 : pht_33; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_450 = 6'h22 == io_execute_update_pht_index ? _pht_T_2 : pht_34; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_451 = 6'h23 == io_execute_update_pht_index ? _pht_T_2 : pht_35; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_452 = 6'h24 == io_execute_update_pht_index ? _pht_T_2 : pht_36; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_453 = 6'h25 == io_execute_update_pht_index ? _pht_T_2 : pht_37; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_454 = 6'h26 == io_execute_update_pht_index ? _pht_T_2 : pht_38; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_455 = 6'h27 == io_execute_update_pht_index ? _pht_T_2 : pht_39; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_456 = 6'h28 == io_execute_update_pht_index ? _pht_T_2 : pht_40; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_457 = 6'h29 == io_execute_update_pht_index ? _pht_T_2 : pht_41; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_458 = 6'h2a == io_execute_update_pht_index ? _pht_T_2 : pht_42; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_459 = 6'h2b == io_execute_update_pht_index ? _pht_T_2 : pht_43; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_460 = 6'h2c == io_execute_update_pht_index ? _pht_T_2 : pht_44; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_461 = 6'h2d == io_execute_update_pht_index ? _pht_T_2 : pht_45; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_462 = 6'h2e == io_execute_update_pht_index ? _pht_T_2 : pht_46; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_463 = 6'h2f == io_execute_update_pht_index ? _pht_T_2 : pht_47; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_464 = 6'h30 == io_execute_update_pht_index ? _pht_T_2 : pht_48; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_465 = 6'h31 == io_execute_update_pht_index ? _pht_T_2 : pht_49; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_466 = 6'h32 == io_execute_update_pht_index ? _pht_T_2 : pht_50; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_467 = 6'h33 == io_execute_update_pht_index ? _pht_T_2 : pht_51; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_468 = 6'h34 == io_execute_update_pht_index ? _pht_T_2 : pht_52; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_469 = 6'h35 == io_execute_update_pht_index ? _pht_T_2 : pht_53; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_470 = 6'h36 == io_execute_update_pht_index ? _pht_T_2 : pht_54; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_471 = 6'h37 == io_execute_update_pht_index ? _pht_T_2 : pht_55; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_472 = 6'h38 == io_execute_update_pht_index ? _pht_T_2 : pht_56; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_473 = 6'h39 == io_execute_update_pht_index ? _pht_T_2 : pht_57; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_474 = 6'h3a == io_execute_update_pht_index ? _pht_T_2 : pht_58; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_475 = 6'h3b == io_execute_update_pht_index ? _pht_T_2 : pht_59; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_476 = 6'h3c == io_execute_update_pht_index ? _pht_T_2 : pht_60; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_477 = 6'h3d == io_execute_update_pht_index ? _pht_T_2 : pht_61; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_478 = 6'h3e == io_execute_update_pht_index ? _pht_T_2 : pht_62; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _GEN_479 = 6'h3f == io_execute_update_pht_index ? _pht_T_2 : pht_63; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 142:{31,31}]
  wire [1:0] _pht_T_3 = io_execute_branch ? 2'h3 : 2'h2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 145:37]
  wire [1:0] _GEN_480 = 6'h0 == io_execute_update_pht_index ? _pht_T_3 : pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_481 = 6'h1 == io_execute_update_pht_index ? _pht_T_3 : pht_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_482 = 6'h2 == io_execute_update_pht_index ? _pht_T_3 : pht_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_483 = 6'h3 == io_execute_update_pht_index ? _pht_T_3 : pht_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_484 = 6'h4 == io_execute_update_pht_index ? _pht_T_3 : pht_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_485 = 6'h5 == io_execute_update_pht_index ? _pht_T_3 : pht_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_486 = 6'h6 == io_execute_update_pht_index ? _pht_T_3 : pht_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_487 = 6'h7 == io_execute_update_pht_index ? _pht_T_3 : pht_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_488 = 6'h8 == io_execute_update_pht_index ? _pht_T_3 : pht_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_489 = 6'h9 == io_execute_update_pht_index ? _pht_T_3 : pht_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_490 = 6'ha == io_execute_update_pht_index ? _pht_T_3 : pht_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_491 = 6'hb == io_execute_update_pht_index ? _pht_T_3 : pht_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_492 = 6'hc == io_execute_update_pht_index ? _pht_T_3 : pht_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_493 = 6'hd == io_execute_update_pht_index ? _pht_T_3 : pht_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_494 = 6'he == io_execute_update_pht_index ? _pht_T_3 : pht_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_495 = 6'hf == io_execute_update_pht_index ? _pht_T_3 : pht_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_496 = 6'h10 == io_execute_update_pht_index ? _pht_T_3 : pht_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_497 = 6'h11 == io_execute_update_pht_index ? _pht_T_3 : pht_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_498 = 6'h12 == io_execute_update_pht_index ? _pht_T_3 : pht_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_499 = 6'h13 == io_execute_update_pht_index ? _pht_T_3 : pht_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_500 = 6'h14 == io_execute_update_pht_index ? _pht_T_3 : pht_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_501 = 6'h15 == io_execute_update_pht_index ? _pht_T_3 : pht_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_502 = 6'h16 == io_execute_update_pht_index ? _pht_T_3 : pht_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_503 = 6'h17 == io_execute_update_pht_index ? _pht_T_3 : pht_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_504 = 6'h18 == io_execute_update_pht_index ? _pht_T_3 : pht_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_505 = 6'h19 == io_execute_update_pht_index ? _pht_T_3 : pht_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_506 = 6'h1a == io_execute_update_pht_index ? _pht_T_3 : pht_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_507 = 6'h1b == io_execute_update_pht_index ? _pht_T_3 : pht_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_508 = 6'h1c == io_execute_update_pht_index ? _pht_T_3 : pht_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_509 = 6'h1d == io_execute_update_pht_index ? _pht_T_3 : pht_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_510 = 6'h1e == io_execute_update_pht_index ? _pht_T_3 : pht_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_511 = 6'h1f == io_execute_update_pht_index ? _pht_T_3 : pht_31; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_512 = 6'h20 == io_execute_update_pht_index ? _pht_T_3 : pht_32; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_513 = 6'h21 == io_execute_update_pht_index ? _pht_T_3 : pht_33; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_514 = 6'h22 == io_execute_update_pht_index ? _pht_T_3 : pht_34; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_515 = 6'h23 == io_execute_update_pht_index ? _pht_T_3 : pht_35; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_516 = 6'h24 == io_execute_update_pht_index ? _pht_T_3 : pht_36; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_517 = 6'h25 == io_execute_update_pht_index ? _pht_T_3 : pht_37; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_518 = 6'h26 == io_execute_update_pht_index ? _pht_T_3 : pht_38; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_519 = 6'h27 == io_execute_update_pht_index ? _pht_T_3 : pht_39; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_520 = 6'h28 == io_execute_update_pht_index ? _pht_T_3 : pht_40; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_521 = 6'h29 == io_execute_update_pht_index ? _pht_T_3 : pht_41; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_522 = 6'h2a == io_execute_update_pht_index ? _pht_T_3 : pht_42; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_523 = 6'h2b == io_execute_update_pht_index ? _pht_T_3 : pht_43; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_524 = 6'h2c == io_execute_update_pht_index ? _pht_T_3 : pht_44; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_525 = 6'h2d == io_execute_update_pht_index ? _pht_T_3 : pht_45; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_526 = 6'h2e == io_execute_update_pht_index ? _pht_T_3 : pht_46; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_527 = 6'h2f == io_execute_update_pht_index ? _pht_T_3 : pht_47; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_528 = 6'h30 == io_execute_update_pht_index ? _pht_T_3 : pht_48; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_529 = 6'h31 == io_execute_update_pht_index ? _pht_T_3 : pht_49; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_530 = 6'h32 == io_execute_update_pht_index ? _pht_T_3 : pht_50; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_531 = 6'h33 == io_execute_update_pht_index ? _pht_T_3 : pht_51; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_532 = 6'h34 == io_execute_update_pht_index ? _pht_T_3 : pht_52; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_533 = 6'h35 == io_execute_update_pht_index ? _pht_T_3 : pht_53; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_534 = 6'h36 == io_execute_update_pht_index ? _pht_T_3 : pht_54; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_535 = 6'h37 == io_execute_update_pht_index ? _pht_T_3 : pht_55; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_536 = 6'h38 == io_execute_update_pht_index ? _pht_T_3 : pht_56; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_537 = 6'h39 == io_execute_update_pht_index ? _pht_T_3 : pht_57; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_538 = 6'h3a == io_execute_update_pht_index ? _pht_T_3 : pht_58; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_539 = 6'h3b == io_execute_update_pht_index ? _pht_T_3 : pht_59; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_540 = 6'h3c == io_execute_update_pht_index ? _pht_T_3 : pht_60; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_541 = 6'h3d == io_execute_update_pht_index ? _pht_T_3 : pht_61; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_542 = 6'h3e == io_execute_update_pht_index ? _pht_T_3 : pht_62; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_543 = 6'h3f == io_execute_update_pht_index ? _pht_T_3 : pht_63; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 145:{31,31}]
  wire [1:0] _GEN_544 = 2'h3 == _GEN_287 ? _GEN_480 : pht_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_545 = 2'h3 == _GEN_287 ? _GEN_481 : pht_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_546 = 2'h3 == _GEN_287 ? _GEN_482 : pht_2; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_547 = 2'h3 == _GEN_287 ? _GEN_483 : pht_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_548 = 2'h3 == _GEN_287 ? _GEN_484 : pht_4; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_549 = 2'h3 == _GEN_287 ? _GEN_485 : pht_5; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_550 = 2'h3 == _GEN_287 ? _GEN_486 : pht_6; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_551 = 2'h3 == _GEN_287 ? _GEN_487 : pht_7; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_552 = 2'h3 == _GEN_287 ? _GEN_488 : pht_8; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_553 = 2'h3 == _GEN_287 ? _GEN_489 : pht_9; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_554 = 2'h3 == _GEN_287 ? _GEN_490 : pht_10; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_555 = 2'h3 == _GEN_287 ? _GEN_491 : pht_11; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_556 = 2'h3 == _GEN_287 ? _GEN_492 : pht_12; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_557 = 2'h3 == _GEN_287 ? _GEN_493 : pht_13; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_558 = 2'h3 == _GEN_287 ? _GEN_494 : pht_14; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_559 = 2'h3 == _GEN_287 ? _GEN_495 : pht_15; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_560 = 2'h3 == _GEN_287 ? _GEN_496 : pht_16; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_561 = 2'h3 == _GEN_287 ? _GEN_497 : pht_17; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_562 = 2'h3 == _GEN_287 ? _GEN_498 : pht_18; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_563 = 2'h3 == _GEN_287 ? _GEN_499 : pht_19; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_564 = 2'h3 == _GEN_287 ? _GEN_500 : pht_20; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_565 = 2'h3 == _GEN_287 ? _GEN_501 : pht_21; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_566 = 2'h3 == _GEN_287 ? _GEN_502 : pht_22; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_567 = 2'h3 == _GEN_287 ? _GEN_503 : pht_23; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_568 = 2'h3 == _GEN_287 ? _GEN_504 : pht_24; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_569 = 2'h3 == _GEN_287 ? _GEN_505 : pht_25; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_570 = 2'h3 == _GEN_287 ? _GEN_506 : pht_26; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_571 = 2'h3 == _GEN_287 ? _GEN_507 : pht_27; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_572 = 2'h3 == _GEN_287 ? _GEN_508 : pht_28; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_573 = 2'h3 == _GEN_287 ? _GEN_509 : pht_29; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_574 = 2'h3 == _GEN_287 ? _GEN_510 : pht_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_575 = 2'h3 == _GEN_287 ? _GEN_511 : pht_31; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_576 = 2'h3 == _GEN_287 ? _GEN_512 : pht_32; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_577 = 2'h3 == _GEN_287 ? _GEN_513 : pht_33; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_578 = 2'h3 == _GEN_287 ? _GEN_514 : pht_34; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_579 = 2'h3 == _GEN_287 ? _GEN_515 : pht_35; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_580 = 2'h3 == _GEN_287 ? _GEN_516 : pht_36; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_581 = 2'h3 == _GEN_287 ? _GEN_517 : pht_37; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_582 = 2'h3 == _GEN_287 ? _GEN_518 : pht_38; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_583 = 2'h3 == _GEN_287 ? _GEN_519 : pht_39; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_584 = 2'h3 == _GEN_287 ? _GEN_520 : pht_40; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_585 = 2'h3 == _GEN_287 ? _GEN_521 : pht_41; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_586 = 2'h3 == _GEN_287 ? _GEN_522 : pht_42; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_587 = 2'h3 == _GEN_287 ? _GEN_523 : pht_43; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_588 = 2'h3 == _GEN_287 ? _GEN_524 : pht_44; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_589 = 2'h3 == _GEN_287 ? _GEN_525 : pht_45; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_590 = 2'h3 == _GEN_287 ? _GEN_526 : pht_46; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_591 = 2'h3 == _GEN_287 ? _GEN_527 : pht_47; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_592 = 2'h3 == _GEN_287 ? _GEN_528 : pht_48; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_593 = 2'h3 == _GEN_287 ? _GEN_529 : pht_49; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_594 = 2'h3 == _GEN_287 ? _GEN_530 : pht_50; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_595 = 2'h3 == _GEN_287 ? _GEN_531 : pht_51; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_596 = 2'h3 == _GEN_287 ? _GEN_532 : pht_52; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_597 = 2'h3 == _GEN_287 ? _GEN_533 : pht_53; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_598 = 2'h3 == _GEN_287 ? _GEN_534 : pht_54; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_599 = 2'h3 == _GEN_287 ? _GEN_535 : pht_55; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_600 = 2'h3 == _GEN_287 ? _GEN_536 : pht_56; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_601 = 2'h3 == _GEN_287 ? _GEN_537 : pht_57; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_602 = 2'h3 == _GEN_287 ? _GEN_538 : pht_58; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_603 = 2'h3 == _GEN_287 ? _GEN_539 : pht_59; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_604 = 2'h3 == _GEN_287 ? _GEN_540 : pht_60; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_605 = 2'h3 == _GEN_287 ? _GEN_541 : pht_61; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_606 = 2'h3 == _GEN_287 ? _GEN_542 : pht_62; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_607 = 2'h3 == _GEN_287 ? _GEN_543 : pht_63; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26 134:35]
  wire [1:0] _GEN_608 = 2'h2 == _GEN_287 ? _GEN_416 : _GEN_544; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_609 = 2'h2 == _GEN_287 ? _GEN_417 : _GEN_545; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_610 = 2'h2 == _GEN_287 ? _GEN_418 : _GEN_546; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_611 = 2'h2 == _GEN_287 ? _GEN_419 : _GEN_547; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_612 = 2'h2 == _GEN_287 ? _GEN_420 : _GEN_548; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_613 = 2'h2 == _GEN_287 ? _GEN_421 : _GEN_549; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_614 = 2'h2 == _GEN_287 ? _GEN_422 : _GEN_550; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_615 = 2'h2 == _GEN_287 ? _GEN_423 : _GEN_551; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_616 = 2'h2 == _GEN_287 ? _GEN_424 : _GEN_552; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_617 = 2'h2 == _GEN_287 ? _GEN_425 : _GEN_553; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_618 = 2'h2 == _GEN_287 ? _GEN_426 : _GEN_554; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_619 = 2'h2 == _GEN_287 ? _GEN_427 : _GEN_555; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_620 = 2'h2 == _GEN_287 ? _GEN_428 : _GEN_556; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_621 = 2'h2 == _GEN_287 ? _GEN_429 : _GEN_557; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_622 = 2'h2 == _GEN_287 ? _GEN_430 : _GEN_558; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_623 = 2'h2 == _GEN_287 ? _GEN_431 : _GEN_559; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_624 = 2'h2 == _GEN_287 ? _GEN_432 : _GEN_560; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_625 = 2'h2 == _GEN_287 ? _GEN_433 : _GEN_561; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_626 = 2'h2 == _GEN_287 ? _GEN_434 : _GEN_562; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_627 = 2'h2 == _GEN_287 ? _GEN_435 : _GEN_563; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_628 = 2'h2 == _GEN_287 ? _GEN_436 : _GEN_564; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_629 = 2'h2 == _GEN_287 ? _GEN_437 : _GEN_565; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_630 = 2'h2 == _GEN_287 ? _GEN_438 : _GEN_566; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_631 = 2'h2 == _GEN_287 ? _GEN_439 : _GEN_567; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_632 = 2'h2 == _GEN_287 ? _GEN_440 : _GEN_568; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_633 = 2'h2 == _GEN_287 ? _GEN_441 : _GEN_569; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_634 = 2'h2 == _GEN_287 ? _GEN_442 : _GEN_570; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_635 = 2'h2 == _GEN_287 ? _GEN_443 : _GEN_571; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_636 = 2'h2 == _GEN_287 ? _GEN_444 : _GEN_572; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_637 = 2'h2 == _GEN_287 ? _GEN_445 : _GEN_573; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_638 = 2'h2 == _GEN_287 ? _GEN_446 : _GEN_574; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_639 = 2'h2 == _GEN_287 ? _GEN_447 : _GEN_575; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_640 = 2'h2 == _GEN_287 ? _GEN_448 : _GEN_576; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_641 = 2'h2 == _GEN_287 ? _GEN_449 : _GEN_577; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_642 = 2'h2 == _GEN_287 ? _GEN_450 : _GEN_578; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_643 = 2'h2 == _GEN_287 ? _GEN_451 : _GEN_579; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_644 = 2'h2 == _GEN_287 ? _GEN_452 : _GEN_580; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_645 = 2'h2 == _GEN_287 ? _GEN_453 : _GEN_581; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_646 = 2'h2 == _GEN_287 ? _GEN_454 : _GEN_582; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_647 = 2'h2 == _GEN_287 ? _GEN_455 : _GEN_583; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_648 = 2'h2 == _GEN_287 ? _GEN_456 : _GEN_584; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_649 = 2'h2 == _GEN_287 ? _GEN_457 : _GEN_585; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_650 = 2'h2 == _GEN_287 ? _GEN_458 : _GEN_586; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_651 = 2'h2 == _GEN_287 ? _GEN_459 : _GEN_587; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_652 = 2'h2 == _GEN_287 ? _GEN_460 : _GEN_588; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_653 = 2'h2 == _GEN_287 ? _GEN_461 : _GEN_589; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_654 = 2'h2 == _GEN_287 ? _GEN_462 : _GEN_590; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_655 = 2'h2 == _GEN_287 ? _GEN_463 : _GEN_591; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_656 = 2'h2 == _GEN_287 ? _GEN_464 : _GEN_592; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_657 = 2'h2 == _GEN_287 ? _GEN_465 : _GEN_593; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_658 = 2'h2 == _GEN_287 ? _GEN_466 : _GEN_594; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_659 = 2'h2 == _GEN_287 ? _GEN_467 : _GEN_595; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_660 = 2'h2 == _GEN_287 ? _GEN_468 : _GEN_596; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_661 = 2'h2 == _GEN_287 ? _GEN_469 : _GEN_597; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_662 = 2'h2 == _GEN_287 ? _GEN_470 : _GEN_598; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_663 = 2'h2 == _GEN_287 ? _GEN_471 : _GEN_599; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_664 = 2'h2 == _GEN_287 ? _GEN_472 : _GEN_600; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_665 = 2'h2 == _GEN_287 ? _GEN_473 : _GEN_601; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_666 = 2'h2 == _GEN_287 ? _GEN_474 : _GEN_602; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_667 = 2'h2 == _GEN_287 ? _GEN_475 : _GEN_603; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_668 = 2'h2 == _GEN_287 ? _GEN_476 : _GEN_604; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_669 = 2'h2 == _GEN_287 ? _GEN_477 : _GEN_605; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_670 = 2'h2 == _GEN_287 ? _GEN_478 : _GEN_606; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  wire [1:0] _GEN_671 = 2'h2 == _GEN_287 ? _GEN_479 : _GEN_607; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
  assign io_decode_branch_inst = _io_decode_branch_inst_T_1 & _io_decode_branch_inst_T_3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 114:41]
  assign io_decode_branch = io_decode_branch_inst & (_GEN_127 == 2'h2 | _GEN_127 == 2'h3); // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 126:27]
  assign io_decode_target = io_decode_pc + io_decode_info_imm; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 115:36]
  assign io_decode_update_pht_index = 5'h1f == io_decode_pc[6:2] ? bht_31 : _GEN_158; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 127:{30,30}]
  assign io_instBuffer_pht_index_0 = 5'h1f == io_instBuffer_pc_0[6:2] ? bht_31 : _GEN_30; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  assign io_instBuffer_pht_index_1 = 5'h1f == io_instBuffer_pc_1[6:2] ? bht_31 : _GEN_62; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 122:{32,32}]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_0 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h0 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_0 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_1 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_1 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_2 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h2 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_2 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_3 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h3 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_3 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_4 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h4 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_4 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_5 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h5 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_5 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_6 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h6 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_6 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_7 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h7 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_7 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_8 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h8 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_8 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_9 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h9 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_9 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_10 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'ha == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_10 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_11 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'hb == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_11 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_12 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'hc == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_12 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_13 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'hd == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_13 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_14 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'he == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_14 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_15 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'hf == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_15 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_16 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h10 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_16 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_17 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h11 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_17 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_18 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h12 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_18 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_19 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h13 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_19 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_20 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h14 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_20 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_21 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h15 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_21 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_22 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h16 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_22 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_23 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h17 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_23 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_24 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h18 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_24 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_25 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h19 == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_25 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_26 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1a == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_26 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_27 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1b == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_27 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_28 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1c == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_28 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_29 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1d == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_29 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_30 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1e == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_30 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
      bht_31 <= 6'h0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 117:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (5'h1f == update_bht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
        bht_31 <= _bht_T_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 133:27]
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_0 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h0 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_0 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_0 <= _GEN_352;
      end else begin
        pht_0 <= _GEN_608;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_1 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_1 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_1 <= _GEN_353;
      end else begin
        pht_1 <= _GEN_609;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_2 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_2 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_2 <= _GEN_354;
      end else begin
        pht_2 <= _GEN_610;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_3 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_3 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_3 <= _GEN_355;
      end else begin
        pht_3 <= _GEN_611;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_4 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h4 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_4 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_4 <= _GEN_356;
      end else begin
        pht_4 <= _GEN_612;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_5 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h5 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_5 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_5 <= _GEN_357;
      end else begin
        pht_5 <= _GEN_613;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_6 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h6 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_6 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_6 <= _GEN_358;
      end else begin
        pht_6 <= _GEN_614;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_7 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h7 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_7 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_7 <= _GEN_359;
      end else begin
        pht_7 <= _GEN_615;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_8 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h8 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_8 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_8 <= _GEN_360;
      end else begin
        pht_8 <= _GEN_616;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_9 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h9 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_9 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_9 <= _GEN_361;
      end else begin
        pht_9 <= _GEN_617;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_10 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'ha == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_10 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_10 <= _GEN_362;
      end else begin
        pht_10 <= _GEN_618;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_11 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'hb == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_11 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_11 <= _GEN_363;
      end else begin
        pht_11 <= _GEN_619;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_12 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'hc == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_12 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_12 <= _GEN_364;
      end else begin
        pht_12 <= _GEN_620;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_13 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'hd == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_13 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_13 <= _GEN_365;
      end else begin
        pht_13 <= _GEN_621;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_14 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'he == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_14 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_14 <= _GEN_366;
      end else begin
        pht_14 <= _GEN_622;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_15 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'hf == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_15 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_15 <= _GEN_367;
      end else begin
        pht_15 <= _GEN_623;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_16 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h10 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_16 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_16 <= _GEN_368;
      end else begin
        pht_16 <= _GEN_624;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_17 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h11 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_17 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_17 <= _GEN_369;
      end else begin
        pht_17 <= _GEN_625;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_18 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h12 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_18 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_18 <= _GEN_370;
      end else begin
        pht_18 <= _GEN_626;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_19 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h13 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_19 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_19 <= _GEN_371;
      end else begin
        pht_19 <= _GEN_627;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_20 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h14 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_20 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_20 <= _GEN_372;
      end else begin
        pht_20 <= _GEN_628;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_21 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h15 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_21 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_21 <= _GEN_373;
      end else begin
        pht_21 <= _GEN_629;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_22 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h16 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_22 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_22 <= _GEN_374;
      end else begin
        pht_22 <= _GEN_630;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_23 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h17 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_23 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_23 <= _GEN_375;
      end else begin
        pht_23 <= _GEN_631;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_24 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h18 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_24 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_24 <= _GEN_376;
      end else begin
        pht_24 <= _GEN_632;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_25 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h19 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_25 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_25 <= _GEN_377;
      end else begin
        pht_25 <= _GEN_633;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_26 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1a == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_26 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_26 <= _GEN_378;
      end else begin
        pht_26 <= _GEN_634;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_27 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1b == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_27 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_27 <= _GEN_379;
      end else begin
        pht_27 <= _GEN_635;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_28 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1c == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_28 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_28 <= _GEN_380;
      end else begin
        pht_28 <= _GEN_636;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_29 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1d == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_29 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_29 <= _GEN_381;
      end else begin
        pht_29 <= _GEN_637;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_30 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1e == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_30 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_30 <= _GEN_382;
      end else begin
        pht_30 <= _GEN_638;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_31 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h1f == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_31 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_31 <= _GEN_383;
      end else begin
        pht_31 <= _GEN_639;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_32 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h20 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_32 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_32 <= _GEN_384;
      end else begin
        pht_32 <= _GEN_640;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_33 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h21 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_33 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_33 <= _GEN_385;
      end else begin
        pht_33 <= _GEN_641;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_34 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h22 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_34 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_34 <= _GEN_386;
      end else begin
        pht_34 <= _GEN_642;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_35 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h23 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_35 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_35 <= _GEN_387;
      end else begin
        pht_35 <= _GEN_643;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_36 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h24 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_36 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_36 <= _GEN_388;
      end else begin
        pht_36 <= _GEN_644;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_37 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h25 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_37 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_37 <= _GEN_389;
      end else begin
        pht_37 <= _GEN_645;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_38 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h26 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_38 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_38 <= _GEN_390;
      end else begin
        pht_38 <= _GEN_646;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_39 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h27 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_39 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_39 <= _GEN_391;
      end else begin
        pht_39 <= _GEN_647;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_40 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h28 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_40 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_40 <= _GEN_392;
      end else begin
        pht_40 <= _GEN_648;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_41 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h29 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_41 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_41 <= _GEN_393;
      end else begin
        pht_41 <= _GEN_649;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_42 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2a == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_42 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_42 <= _GEN_394;
      end else begin
        pht_42 <= _GEN_650;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_43 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2b == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_43 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_43 <= _GEN_395;
      end else begin
        pht_43 <= _GEN_651;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_44 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2c == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_44 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_44 <= _GEN_396;
      end else begin
        pht_44 <= _GEN_652;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_45 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2d == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_45 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_45 <= _GEN_397;
      end else begin
        pht_45 <= _GEN_653;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_46 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2e == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_46 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_46 <= _GEN_398;
      end else begin
        pht_46 <= _GEN_654;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_47 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h2f == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_47 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_47 <= _GEN_399;
      end else begin
        pht_47 <= _GEN_655;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_48 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h30 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_48 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_48 <= _GEN_400;
      end else begin
        pht_48 <= _GEN_656;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_49 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h31 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_49 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_49 <= _GEN_401;
      end else begin
        pht_49 <= _GEN_657;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_50 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h32 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_50 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_50 <= _GEN_402;
      end else begin
        pht_50 <= _GEN_658;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_51 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h33 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_51 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_51 <= _GEN_403;
      end else begin
        pht_51 <= _GEN_659;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_52 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h34 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_52 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_52 <= _GEN_404;
      end else begin
        pht_52 <= _GEN_660;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_53 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h35 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_53 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_53 <= _GEN_405;
      end else begin
        pht_53 <= _GEN_661;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_54 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h36 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_54 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_54 <= _GEN_406;
      end else begin
        pht_54 <= _GEN_662;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_55 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h37 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_55 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_55 <= _GEN_407;
      end else begin
        pht_55 <= _GEN_663;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_56 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h38 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_56 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_56 <= _GEN_408;
      end else begin
        pht_56 <= _GEN_664;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_57 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h39 == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_57 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_57 <= _GEN_409;
      end else begin
        pht_57 <= _GEN_665;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_58 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3a == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_58 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_58 <= _GEN_410;
      end else begin
        pht_58 <= _GEN_666;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_59 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3b == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_59 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_59 <= _GEN_411;
      end else begin
        pht_59 <= _GEN_667;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_60 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3c == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_60 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_60 <= _GEN_412;
      end else begin
        pht_60 <= _GEN_668;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_61 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3d == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_61 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_61 <= _GEN_413;
      end else begin
        pht_61 <= _GEN_669;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_62 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3e == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_62 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_62 <= _GEN_414;
      end else begin
        pht_62 <= _GEN_670;
      end
    end
    if (reset) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
      pht_63 <= 2'h3; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 118:26]
    end else if (io_execute_branch_inst) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 132:32]
      if (2'h0 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        if (6'h3f == io_execute_update_pht_index) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
          pht_63 <= _pht_T; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 136:31]
        end
      end else if (2'h1 == _GEN_287) begin // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 134:35]
        pht_63 <= _GEN_415;
      end else begin
        pht_63 <= _GEN_671;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bht_0 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  bht_1 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  bht_2 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  bht_3 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  bht_4 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  bht_5 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  bht_6 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  bht_7 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  bht_8 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  bht_9 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  bht_10 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  bht_11 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  bht_12 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  bht_13 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  bht_14 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  bht_15 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  bht_16 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  bht_17 = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  bht_18 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  bht_19 = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  bht_20 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  bht_21 = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  bht_22 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  bht_23 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  bht_24 = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  bht_25 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  bht_26 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  bht_27 = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  bht_28 = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  bht_29 = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  bht_30 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  bht_31 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  pht_0 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  pht_1 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  pht_2 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  pht_3 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  pht_4 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  pht_5 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  pht_6 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  pht_7 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  pht_8 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  pht_9 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  pht_10 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  pht_11 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  pht_12 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  pht_13 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  pht_14 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  pht_15 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  pht_16 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  pht_17 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  pht_18 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  pht_19 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  pht_20 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  pht_21 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  pht_22 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  pht_23 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  pht_24 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  pht_25 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  pht_26 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  pht_27 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  pht_28 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  pht_29 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  pht_30 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  pht_31 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  pht_32 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pht_33 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pht_34 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pht_35 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pht_36 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pht_37 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pht_38 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pht_39 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pht_40 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pht_41 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pht_42 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pht_43 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pht_44 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pht_45 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pht_46 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pht_47 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  pht_48 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  pht_49 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  pht_50 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  pht_51 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  pht_52 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  pht_53 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  pht_54 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  pht_55 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  pht_56 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  pht_57 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  pht_58 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  pht_59 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  pht_60 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  pht_61 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  pht_62 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  pht_63 = _RAND_95[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BranchPredictorUnit(
  input         clock,
  input         reset,
  input  [63:0] io_decode_pc, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input         io_decode_info_valid, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [2:0]  io_decode_info_fusel, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [6:0]  io_decode_info_op, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [63:0] io_decode_info_imm, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [5:0]  io_decode_pht_index, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  output        io_decode_branch_inst, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  output        io_decode_branch, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  output [63:0] io_decode_target, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  output [5:0]  io_decode_update_pht_index, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [63:0] io_instBuffer_pc_0, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [63:0] io_instBuffer_pc_1, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  output [5:0]  io_instBuffer_pht_index_0, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  output [5:0]  io_instBuffer_pht_index_1, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [63:0] io_execute_pc, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input  [5:0]  io_execute_update_pht_index, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input         io_execute_branch_inst, // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
  input         io_execute_branch // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 36:14]
);
  wire  adaptive_predictor_clock; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire  adaptive_predictor_reset; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [63:0] adaptive_predictor_io_decode_pc; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire  adaptive_predictor_io_decode_info_valid; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [2:0] adaptive_predictor_io_decode_info_fusel; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [6:0] adaptive_predictor_io_decode_info_op; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [63:0] adaptive_predictor_io_decode_info_imm; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [5:0] adaptive_predictor_io_decode_pht_index; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire  adaptive_predictor_io_decode_branch_inst; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire  adaptive_predictor_io_decode_branch; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [63:0] adaptive_predictor_io_decode_target; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [5:0] adaptive_predictor_io_decode_update_pht_index; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [63:0] adaptive_predictor_io_instBuffer_pc_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [63:0] adaptive_predictor_io_instBuffer_pc_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [5:0] adaptive_predictor_io_instBuffer_pht_index_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [5:0] adaptive_predictor_io_instBuffer_pht_index_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [63:0] adaptive_predictor_io_execute_pc; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire [5:0] adaptive_predictor_io_execute_update_pht_index; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire  adaptive_predictor_io_execute_branch_inst; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  wire  adaptive_predictor_io_execute_branch; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
  AdaptiveTwoLevelPredictor adaptive_predictor ( // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 39:36]
    .clock(adaptive_predictor_clock),
    .reset(adaptive_predictor_reset),
    .io_decode_pc(adaptive_predictor_io_decode_pc),
    .io_decode_info_valid(adaptive_predictor_io_decode_info_valid),
    .io_decode_info_fusel(adaptive_predictor_io_decode_info_fusel),
    .io_decode_info_op(adaptive_predictor_io_decode_info_op),
    .io_decode_info_imm(adaptive_predictor_io_decode_info_imm),
    .io_decode_pht_index(adaptive_predictor_io_decode_pht_index),
    .io_decode_branch_inst(adaptive_predictor_io_decode_branch_inst),
    .io_decode_branch(adaptive_predictor_io_decode_branch),
    .io_decode_target(adaptive_predictor_io_decode_target),
    .io_decode_update_pht_index(adaptive_predictor_io_decode_update_pht_index),
    .io_instBuffer_pc_0(adaptive_predictor_io_instBuffer_pc_0),
    .io_instBuffer_pc_1(adaptive_predictor_io_instBuffer_pc_1),
    .io_instBuffer_pht_index_0(adaptive_predictor_io_instBuffer_pht_index_0),
    .io_instBuffer_pht_index_1(adaptive_predictor_io_instBuffer_pht_index_1),
    .io_execute_pc(adaptive_predictor_io_execute_pc),
    .io_execute_update_pht_index(adaptive_predictor_io_execute_update_pht_index),
    .io_execute_branch_inst(adaptive_predictor_io_execute_branch_inst),
    .io_execute_branch(adaptive_predictor_io_execute_branch)
  );
  assign io_decode_branch_inst = adaptive_predictor_io_decode_branch_inst; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign io_decode_branch = adaptive_predictor_io_decode_branch; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign io_decode_target = adaptive_predictor_io_decode_target; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign io_decode_update_pht_index = adaptive_predictor_io_decode_update_pht_index; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign io_instBuffer_pht_index_0 = adaptive_predictor_io_instBuffer_pht_index_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign io_instBuffer_pht_index_1 = adaptive_predictor_io_instBuffer_pht_index_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_clock = clock;
  assign adaptive_predictor_reset = reset;
  assign adaptive_predictor_io_decode_pc = io_decode_pc; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_decode_info_valid = io_decode_info_valid; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_decode_info_fusel = io_decode_info_fusel; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_decode_info_op = io_decode_info_op; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_decode_info_imm = io_decode_info_imm; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_decode_pht_index = io_decode_pht_index; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_instBuffer_pc_0 = io_instBuffer_pc_0; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_instBuffer_pc_1 = io_instBuffer_pc_1; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_execute_pc = io_execute_pc; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_execute_update_pht_index = io_execute_update_pht_index; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_execute_branch_inst = io_execute_branch_inst; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
  assign adaptive_predictor_io_execute_branch = io_execute_branch; // @[playground/src/pipeline/fetch/BranchPredictorUnit.scala 40:8]
endmodule
module InstFifo(
  input         clock,
  input         reset,
  input         io_do_flush, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_wen_0, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_wen_1, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input  [63:0] io_write_0_inst, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input  [5:0]  io_write_0_pht_index, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_write_0_addr_misaligned, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_write_0_access_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_write_0_page_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input  [63:0] io_write_0_pc, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input  [63:0] io_write_1_inst, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input  [5:0]  io_write_1_pht_index, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_write_1_addr_misaligned, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_write_1_access_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_write_1_page_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input  [63:0] io_write_1_pc, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_full, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_decoderUint_allow_to_go_0, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  input         io_decoderUint_allow_to_go_1, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output [63:0] io_decoderUint_inst_0_inst, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output [5:0]  io_decoderUint_inst_0_pht_index, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_inst_0_addr_misaligned, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_inst_0_access_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_inst_0_page_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output [63:0] io_decoderUint_inst_0_pc, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output [63:0] io_decoderUint_inst_1_inst, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_inst_1_addr_misaligned, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_inst_1_access_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_inst_1_page_fault, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output [63:0] io_decoderUint_inst_1_pc, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_info_empty, // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
  output        io_decoderUint_info_almost_empty // @[playground/src/pipeline/fetch/InstFifo.scala 20:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] buffer_0_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_0_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_0_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_0_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_0_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_0_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_2_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_2_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_2_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_2_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_2_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_2_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_3_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_3_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_3_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_3_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_3_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_3_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_4_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_4_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_4_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_4_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_4_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_4_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_5_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_5_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_5_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_5_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_5_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_5_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_6_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_6_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_6_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_6_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_6_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_6_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_7_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [5:0] buffer_7_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_7_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_7_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg  buffer_7_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [63:0] buffer_7_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
  reg [2:0] enq_ptr; // @[playground/src/pipeline/fetch/InstFifo.scala 33:24]
  reg [2:0] deq_ptr; // @[playground/src/pipeline/fetch/InstFifo.scala 34:24]
  reg [2:0] count; // @[playground/src/pipeline/fetch/InstFifo.scala 35:24]
  wire  empty = count == 3'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 41:28]
  wire  almost_empty = count == 3'h1; // @[playground/src/pipeline/fetch/InstFifo.scala 42:28]
  wire [63:0] _GEN_6 = 3'h1 == deq_ptr ? buffer_1_inst : buffer_0_inst; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_7 = 3'h1 == deq_ptr ? buffer_1_pht_index : buffer_0_pht_index; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_8 = 3'h1 == deq_ptr ? buffer_1_addr_misaligned : buffer_0_addr_misaligned; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_9 = 3'h1 == deq_ptr ? buffer_1_access_fault : buffer_0_access_fault; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_10 = 3'h1 == deq_ptr ? buffer_1_page_fault : buffer_0_page_fault; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_11 = 3'h1 == deq_ptr ? buffer_1_pc : buffer_0_pc; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_12 = 3'h2 == deq_ptr ? buffer_2_inst : _GEN_6; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_13 = 3'h2 == deq_ptr ? buffer_2_pht_index : _GEN_7; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_14 = 3'h2 == deq_ptr ? buffer_2_addr_misaligned : _GEN_8; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_15 = 3'h2 == deq_ptr ? buffer_2_access_fault : _GEN_9; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_16 = 3'h2 == deq_ptr ? buffer_2_page_fault : _GEN_10; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_17 = 3'h2 == deq_ptr ? buffer_2_pc : _GEN_11; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_18 = 3'h3 == deq_ptr ? buffer_3_inst : _GEN_12; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_19 = 3'h3 == deq_ptr ? buffer_3_pht_index : _GEN_13; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_20 = 3'h3 == deq_ptr ? buffer_3_addr_misaligned : _GEN_14; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_21 = 3'h3 == deq_ptr ? buffer_3_access_fault : _GEN_15; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_22 = 3'h3 == deq_ptr ? buffer_3_page_fault : _GEN_16; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_23 = 3'h3 == deq_ptr ? buffer_3_pc : _GEN_17; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_24 = 3'h4 == deq_ptr ? buffer_4_inst : _GEN_18; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_25 = 3'h4 == deq_ptr ? buffer_4_pht_index : _GEN_19; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_26 = 3'h4 == deq_ptr ? buffer_4_addr_misaligned : _GEN_20; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_27 = 3'h4 == deq_ptr ? buffer_4_access_fault : _GEN_21; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_28 = 3'h4 == deq_ptr ? buffer_4_page_fault : _GEN_22; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_29 = 3'h4 == deq_ptr ? buffer_4_pc : _GEN_23; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_30 = 3'h5 == deq_ptr ? buffer_5_inst : _GEN_24; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_31 = 3'h5 == deq_ptr ? buffer_5_pht_index : _GEN_25; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_32 = 3'h5 == deq_ptr ? buffer_5_addr_misaligned : _GEN_26; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_33 = 3'h5 == deq_ptr ? buffer_5_access_fault : _GEN_27; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_34 = 3'h5 == deq_ptr ? buffer_5_page_fault : _GEN_28; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_35 = 3'h5 == deq_ptr ? buffer_5_pc : _GEN_29; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_36 = 3'h6 == deq_ptr ? buffer_6_inst : _GEN_30; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_37 = 3'h6 == deq_ptr ? buffer_6_pht_index : _GEN_31; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_38 = 3'h6 == deq_ptr ? buffer_6_addr_misaligned : _GEN_32; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_39 = 3'h6 == deq_ptr ? buffer_6_access_fault : _GEN_33; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_40 = 3'h6 == deq_ptr ? buffer_6_page_fault : _GEN_34; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_41 = 3'h6 == deq_ptr ? buffer_6_pc : _GEN_35; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_42 = 3'h7 == deq_ptr ? buffer_7_inst : _GEN_36; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [5:0] _GEN_43 = 3'h7 == deq_ptr ? buffer_7_pht_index : _GEN_37; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_44 = 3'h7 == deq_ptr ? buffer_7_addr_misaligned : _GEN_38; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_45 = 3'h7 == deq_ptr ? buffer_7_access_fault : _GEN_39; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_46 = 3'h7 == deq_ptr ? buffer_7_page_fault : _GEN_40; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_47 = 3'h7 == deq_ptr ? buffer_7_pc : _GEN_41; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [2:0] _io_decoderUint_inst_1_T_1 = deq_ptr + 3'h1; // @[playground/src/pipeline/fetch/InstFifo.scala 58:20]
  wire  _io_decoderUint_inst_1_T_2 = empty | almost_empty; // @[playground/src/pipeline/fetch/InstFifo.scala 60:14]
  wire [63:0] _GEN_54 = 3'h1 == _io_decoderUint_inst_1_T_1 ? buffer_1_inst : buffer_0_inst; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_56 = 3'h1 == _io_decoderUint_inst_1_T_1 ? buffer_1_addr_misaligned : buffer_0_addr_misaligned; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_57 = 3'h1 == _io_decoderUint_inst_1_T_1 ? buffer_1_access_fault : buffer_0_access_fault; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_58 = 3'h1 == _io_decoderUint_inst_1_T_1 ? buffer_1_page_fault : buffer_0_page_fault; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_59 = 3'h1 == _io_decoderUint_inst_1_T_1 ? buffer_1_pc : buffer_0_pc; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_60 = 3'h2 == _io_decoderUint_inst_1_T_1 ? buffer_2_inst : _GEN_54; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_62 = 3'h2 == _io_decoderUint_inst_1_T_1 ? buffer_2_addr_misaligned : _GEN_56; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_63 = 3'h2 == _io_decoderUint_inst_1_T_1 ? buffer_2_access_fault : _GEN_57; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_64 = 3'h2 == _io_decoderUint_inst_1_T_1 ? buffer_2_page_fault : _GEN_58; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_65 = 3'h2 == _io_decoderUint_inst_1_T_1 ? buffer_2_pc : _GEN_59; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_66 = 3'h3 == _io_decoderUint_inst_1_T_1 ? buffer_3_inst : _GEN_60; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_68 = 3'h3 == _io_decoderUint_inst_1_T_1 ? buffer_3_addr_misaligned : _GEN_62; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_69 = 3'h3 == _io_decoderUint_inst_1_T_1 ? buffer_3_access_fault : _GEN_63; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_70 = 3'h3 == _io_decoderUint_inst_1_T_1 ? buffer_3_page_fault : _GEN_64; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_71 = 3'h3 == _io_decoderUint_inst_1_T_1 ? buffer_3_pc : _GEN_65; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_72 = 3'h4 == _io_decoderUint_inst_1_T_1 ? buffer_4_inst : _GEN_66; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_74 = 3'h4 == _io_decoderUint_inst_1_T_1 ? buffer_4_addr_misaligned : _GEN_68; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_75 = 3'h4 == _io_decoderUint_inst_1_T_1 ? buffer_4_access_fault : _GEN_69; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_76 = 3'h4 == _io_decoderUint_inst_1_T_1 ? buffer_4_page_fault : _GEN_70; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_77 = 3'h4 == _io_decoderUint_inst_1_T_1 ? buffer_4_pc : _GEN_71; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_78 = 3'h5 == _io_decoderUint_inst_1_T_1 ? buffer_5_inst : _GEN_72; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_80 = 3'h5 == _io_decoderUint_inst_1_T_1 ? buffer_5_addr_misaligned : _GEN_74; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_81 = 3'h5 == _io_decoderUint_inst_1_T_1 ? buffer_5_access_fault : _GEN_75; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_82 = 3'h5 == _io_decoderUint_inst_1_T_1 ? buffer_5_page_fault : _GEN_76; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_83 = 3'h5 == _io_decoderUint_inst_1_T_1 ? buffer_5_pc : _GEN_77; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_84 = 3'h6 == _io_decoderUint_inst_1_T_1 ? buffer_6_inst : _GEN_78; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_86 = 3'h6 == _io_decoderUint_inst_1_T_1 ? buffer_6_addr_misaligned : _GEN_80; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_87 = 3'h6 == _io_decoderUint_inst_1_T_1 ? buffer_6_access_fault : _GEN_81; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_88 = 3'h6 == _io_decoderUint_inst_1_T_1 ? buffer_6_page_fault : _GEN_82; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_89 = 3'h6 == _io_decoderUint_inst_1_T_1 ? buffer_6_pc : _GEN_83; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_90 = 3'h7 == _io_decoderUint_inst_1_T_1 ? buffer_7_inst : _GEN_84; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_92 = 3'h7 == _io_decoderUint_inst_1_T_1 ? buffer_7_addr_misaligned : _GEN_86; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_93 = 3'h7 == _io_decoderUint_inst_1_T_1 ? buffer_7_access_fault : _GEN_87; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire  _GEN_94 = 3'h7 == _io_decoderUint_inst_1_T_1 ? buffer_7_page_fault : _GEN_88; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [63:0] _GEN_95 = 3'h7 == _io_decoderUint_inst_1_T_1 ? buffer_7_pc : _GEN_89; // @[src/main/scala/chisel3/util/Mux.scala 141:{16,16}]
  wire [1:0] _deq_num_T_1 = io_decoderUint_allow_to_go_1 ? 2'h2 : {{1'd0}, io_decoderUint_allow_to_go_0}; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [1:0] deq_num = empty ? 2'h0 : _deq_num_T_1; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [2:0] _GEN_292 = {{1'd0}, deq_num}; // @[playground/src/pipeline/fetch/InstFifo.scala 76:24]
  wire [2:0] _deq_ptr_T_1 = deq_ptr + _GEN_292; // @[playground/src/pipeline/fetch/InstFifo.scala 76:24]
  wire [3:0] _T = {{1'd0}, enq_ptr}; // @[playground/src/pipeline/fetch/InstFifo.scala 84:22]
  wire [63:0] _GEN_97 = 3'h0 == _T[2:0] ? io_write_0_inst : buffer_0_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_98 = 3'h1 == _T[2:0] ? io_write_0_inst : buffer_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_99 = 3'h2 == _T[2:0] ? io_write_0_inst : buffer_2_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_100 = 3'h3 == _T[2:0] ? io_write_0_inst : buffer_3_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_101 = 3'h4 == _T[2:0] ? io_write_0_inst : buffer_4_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_102 = 3'h5 == _T[2:0] ? io_write_0_inst : buffer_5_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_103 = 3'h6 == _T[2:0] ? io_write_0_inst : buffer_6_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_104 = 3'h7 == _T[2:0] ? io_write_0_inst : buffer_7_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_105 = 3'h0 == _T[2:0] ? io_write_0_pht_index : buffer_0_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_106 = 3'h1 == _T[2:0] ? io_write_0_pht_index : buffer_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_107 = 3'h2 == _T[2:0] ? io_write_0_pht_index : buffer_2_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_108 = 3'h3 == _T[2:0] ? io_write_0_pht_index : buffer_3_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_109 = 3'h4 == _T[2:0] ? io_write_0_pht_index : buffer_4_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_110 = 3'h5 == _T[2:0] ? io_write_0_pht_index : buffer_5_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_111 = 3'h6 == _T[2:0] ? io_write_0_pht_index : buffer_6_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [5:0] _GEN_112 = 3'h7 == _T[2:0] ? io_write_0_pht_index : buffer_7_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_113 = 3'h0 == _T[2:0] ? io_write_0_addr_misaligned : buffer_0_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_114 = 3'h1 == _T[2:0] ? io_write_0_addr_misaligned : buffer_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_115 = 3'h2 == _T[2:0] ? io_write_0_addr_misaligned : buffer_2_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_116 = 3'h3 == _T[2:0] ? io_write_0_addr_misaligned : buffer_3_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_117 = 3'h4 == _T[2:0] ? io_write_0_addr_misaligned : buffer_4_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_118 = 3'h5 == _T[2:0] ? io_write_0_addr_misaligned : buffer_5_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_119 = 3'h6 == _T[2:0] ? io_write_0_addr_misaligned : buffer_6_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_120 = 3'h7 == _T[2:0] ? io_write_0_addr_misaligned : buffer_7_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_121 = 3'h0 == _T[2:0] ? io_write_0_access_fault : buffer_0_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_122 = 3'h1 == _T[2:0] ? io_write_0_access_fault : buffer_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_123 = 3'h2 == _T[2:0] ? io_write_0_access_fault : buffer_2_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_124 = 3'h3 == _T[2:0] ? io_write_0_access_fault : buffer_3_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_125 = 3'h4 == _T[2:0] ? io_write_0_access_fault : buffer_4_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_126 = 3'h5 == _T[2:0] ? io_write_0_access_fault : buffer_5_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_127 = 3'h6 == _T[2:0] ? io_write_0_access_fault : buffer_6_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_128 = 3'h7 == _T[2:0] ? io_write_0_access_fault : buffer_7_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_129 = 3'h0 == _T[2:0] ? io_write_0_page_fault : buffer_0_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_130 = 3'h1 == _T[2:0] ? io_write_0_page_fault : buffer_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_131 = 3'h2 == _T[2:0] ? io_write_0_page_fault : buffer_2_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_132 = 3'h3 == _T[2:0] ? io_write_0_page_fault : buffer_3_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_133 = 3'h4 == _T[2:0] ? io_write_0_page_fault : buffer_4_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_134 = 3'h5 == _T[2:0] ? io_write_0_page_fault : buffer_5_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_135 = 3'h6 == _T[2:0] ? io_write_0_page_fault : buffer_6_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire  _GEN_136 = 3'h7 == _T[2:0] ? io_write_0_page_fault : buffer_7_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_137 = 3'h0 == _T[2:0] ? io_write_0_pc : buffer_0_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_138 = 3'h1 == _T[2:0] ? io_write_0_pc : buffer_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_139 = 3'h2 == _T[2:0] ? io_write_0_pc : buffer_2_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_140 = 3'h3 == _T[2:0] ? io_write_0_pc : buffer_3_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_141 = 3'h4 == _T[2:0] ? io_write_0_pc : buffer_4_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_142 = 3'h5 == _T[2:0] ? io_write_0_pc : buffer_5_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_143 = 3'h6 == _T[2:0] ? io_write_0_pc : buffer_6_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_144 = 3'h7 == _T[2:0] ? io_write_0_pc : buffer_7_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23 84:{29,29}]
  wire [63:0] _GEN_145 = io_wen_0 ? _GEN_97 : buffer_0_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_146 = io_wen_0 ? _GEN_98 : buffer_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_147 = io_wen_0 ? _GEN_99 : buffer_2_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_148 = io_wen_0 ? _GEN_100 : buffer_3_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_149 = io_wen_0 ? _GEN_101 : buffer_4_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_150 = io_wen_0 ? _GEN_102 : buffer_5_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_151 = io_wen_0 ? _GEN_103 : buffer_6_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_152 = io_wen_0 ? _GEN_104 : buffer_7_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_153 = io_wen_0 ? _GEN_105 : buffer_0_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_154 = io_wen_0 ? _GEN_106 : buffer_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_155 = io_wen_0 ? _GEN_107 : buffer_2_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_156 = io_wen_0 ? _GEN_108 : buffer_3_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_157 = io_wen_0 ? _GEN_109 : buffer_4_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_158 = io_wen_0 ? _GEN_110 : buffer_5_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_159 = io_wen_0 ? _GEN_111 : buffer_6_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [5:0] _GEN_160 = io_wen_0 ? _GEN_112 : buffer_7_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_161 = io_wen_0 ? _GEN_113 : buffer_0_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_162 = io_wen_0 ? _GEN_114 : buffer_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_163 = io_wen_0 ? _GEN_115 : buffer_2_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_164 = io_wen_0 ? _GEN_116 : buffer_3_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_165 = io_wen_0 ? _GEN_117 : buffer_4_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_166 = io_wen_0 ? _GEN_118 : buffer_5_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_167 = io_wen_0 ? _GEN_119 : buffer_6_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_168 = io_wen_0 ? _GEN_120 : buffer_7_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_169 = io_wen_0 ? _GEN_121 : buffer_0_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_170 = io_wen_0 ? _GEN_122 : buffer_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_171 = io_wen_0 ? _GEN_123 : buffer_2_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_172 = io_wen_0 ? _GEN_124 : buffer_3_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_173 = io_wen_0 ? _GEN_125 : buffer_4_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_174 = io_wen_0 ? _GEN_126 : buffer_5_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_175 = io_wen_0 ? _GEN_127 : buffer_6_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_176 = io_wen_0 ? _GEN_128 : buffer_7_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_177 = io_wen_0 ? _GEN_129 : buffer_0_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_178 = io_wen_0 ? _GEN_130 : buffer_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_179 = io_wen_0 ? _GEN_131 : buffer_2_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_180 = io_wen_0 ? _GEN_132 : buffer_3_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_181 = io_wen_0 ? _GEN_133 : buffer_4_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_182 = io_wen_0 ? _GEN_134 : buffer_5_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_183 = io_wen_0 ? _GEN_135 : buffer_6_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire  _GEN_184 = io_wen_0 ? _GEN_136 : buffer_7_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_185 = io_wen_0 ? _GEN_137 : buffer_0_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_186 = io_wen_0 ? _GEN_138 : buffer_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_187 = io_wen_0 ? _GEN_139 : buffer_2_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_188 = io_wen_0 ? _GEN_140 : buffer_3_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_189 = io_wen_0 ? _GEN_141 : buffer_4_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_190 = io_wen_0 ? _GEN_142 : buffer_5_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_191 = io_wen_0 ? _GEN_143 : buffer_6_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [63:0] _GEN_192 = io_wen_0 ? _GEN_144 : buffer_7_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 83:21 30:23]
  wire [2:0] _T_3 = enq_ptr + 3'h1; // @[playground/src/pipeline/fetch/InstFifo.scala 84:22]
  wire [1:0] enq_num = io_wen_1 ? 2'h2 : {{1'd0}, io_wen_0}; // @[playground/src/pipeline/fetch/InstFifo.scala 96:21 97:15]
  wire [2:0] _GEN_293 = {{1'd0}, enq_num}; // @[playground/src/pipeline/fetch/InstFifo.scala 91:24]
  wire [2:0] _enq_ptr_T_1 = enq_ptr + _GEN_293; // @[playground/src/pipeline/fetch/InstFifo.scala 91:24]
  wire [2:0] _count_T_1 = count + _GEN_293; // @[playground/src/pipeline/fetch/InstFifo.scala 101:40]
  wire [3:0] _GEN_295 = {{1'd0}, _count_T_1}; // @[playground/src/pipeline/fetch/InstFifo.scala 101:50]
  wire [3:0] _count_T_3 = _GEN_295 + 4'h8; // @[playground/src/pipeline/fetch/InstFifo.scala 101:50]
  wire [3:0] _GEN_296 = {{2'd0}, deq_num}; // @[playground/src/pipeline/fetch/InstFifo.scala 101:78]
  wire [3:0] _count_T_5 = _count_T_3 - _GEN_296; // @[playground/src/pipeline/fetch/InstFifo.scala 101:78]
  wire [3:0] _count_T_6 = io_do_flush ? 4'h0 : _count_T_5; // @[playground/src/pipeline/fetch/InstFifo.scala 101:15]
  wire [3:0] _GEN_297 = reset ? 4'h0 : _count_T_6; // @[playground/src/pipeline/fetch/InstFifo.scala 35:{24,24} 101:9]
  assign io_full = count >= 3'h6; // @[playground/src/pipeline/fetch/InstFifo.scala 40:28]
  assign io_decoderUint_inst_0_inst = empty ? 64'h0 : _GEN_42; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_0_pht_index = empty ? 6'h0 : _GEN_43; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_0_addr_misaligned = empty ? 1'h0 : _GEN_44; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_0_access_fault = empty ? 1'h0 : _GEN_45; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_0_page_fault = empty ? 1'h0 : _GEN_46; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_0_pc = empty ? 64'h0 : _GEN_47; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_1_inst = _io_decoderUint_inst_1_T_2 ? 64'h0 : _GEN_90; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_1_addr_misaligned = _io_decoderUint_inst_1_T_2 ? 1'h0 : _GEN_92; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_1_access_fault = _io_decoderUint_inst_1_T_2 ? 1'h0 : _GEN_93; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_1_page_fault = _io_decoderUint_inst_1_T_2 ? 1'h0 : _GEN_94; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_inst_1_pc = _io_decoderUint_inst_1_T_2 ? 64'h0 : _GEN_95; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_decoderUint_info_empty = count == 3'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 41:28]
  assign io_decoderUint_info_almost_empty = count == 3'h1; // @[playground/src/pipeline/fetch/InstFifo.scala 42:28]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_0_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h0 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_0_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_0_inst <= _GEN_145;
      end
    end else begin
      buffer_0_inst <= _GEN_145;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_0_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h0 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_0_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_0_pht_index <= _GEN_153;
      end
    end else begin
      buffer_0_pht_index <= _GEN_153;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_0_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h0 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_0_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_0_addr_misaligned <= _GEN_161;
      end
    end else begin
      buffer_0_addr_misaligned <= _GEN_161;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_0_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h0 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_0_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_0_access_fault <= _GEN_169;
      end
    end else begin
      buffer_0_access_fault <= _GEN_169;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_0_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h0 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_0_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_0_page_fault <= _GEN_177;
      end
    end else begin
      buffer_0_page_fault <= _GEN_177;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_0_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h0 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_0_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_0_pc <= _GEN_185;
      end
    end else begin
      buffer_0_pc <= _GEN_185;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_1_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h1 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_1_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_1_inst <= _GEN_146;
      end
    end else begin
      buffer_1_inst <= _GEN_146;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_1_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h1 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_1_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_1_pht_index <= _GEN_154;
      end
    end else begin
      buffer_1_pht_index <= _GEN_154;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_1_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h1 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_1_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_1_addr_misaligned <= _GEN_162;
      end
    end else begin
      buffer_1_addr_misaligned <= _GEN_162;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_1_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h1 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_1_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_1_access_fault <= _GEN_170;
      end
    end else begin
      buffer_1_access_fault <= _GEN_170;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_1_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h1 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_1_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_1_page_fault <= _GEN_178;
      end
    end else begin
      buffer_1_page_fault <= _GEN_178;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_1_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h1 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_1_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_1_pc <= _GEN_186;
      end
    end else begin
      buffer_1_pc <= _GEN_186;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_2_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h2 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_2_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_2_inst <= _GEN_147;
      end
    end else begin
      buffer_2_inst <= _GEN_147;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_2_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h2 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_2_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_2_pht_index <= _GEN_155;
      end
    end else begin
      buffer_2_pht_index <= _GEN_155;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_2_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h2 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_2_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_2_addr_misaligned <= _GEN_163;
      end
    end else begin
      buffer_2_addr_misaligned <= _GEN_163;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_2_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h2 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_2_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_2_access_fault <= _GEN_171;
      end
    end else begin
      buffer_2_access_fault <= _GEN_171;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_2_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h2 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_2_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_2_page_fault <= _GEN_179;
      end
    end else begin
      buffer_2_page_fault <= _GEN_179;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_2_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h2 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_2_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_2_pc <= _GEN_187;
      end
    end else begin
      buffer_2_pc <= _GEN_187;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_3_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h3 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_3_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_3_inst <= _GEN_148;
      end
    end else begin
      buffer_3_inst <= _GEN_148;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_3_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h3 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_3_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_3_pht_index <= _GEN_156;
      end
    end else begin
      buffer_3_pht_index <= _GEN_156;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_3_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h3 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_3_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_3_addr_misaligned <= _GEN_164;
      end
    end else begin
      buffer_3_addr_misaligned <= _GEN_164;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_3_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h3 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_3_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_3_access_fault <= _GEN_172;
      end
    end else begin
      buffer_3_access_fault <= _GEN_172;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_3_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h3 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_3_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_3_page_fault <= _GEN_180;
      end
    end else begin
      buffer_3_page_fault <= _GEN_180;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_3_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h3 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_3_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_3_pc <= _GEN_188;
      end
    end else begin
      buffer_3_pc <= _GEN_188;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_4_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h4 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_4_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_4_inst <= _GEN_149;
      end
    end else begin
      buffer_4_inst <= _GEN_149;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_4_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h4 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_4_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_4_pht_index <= _GEN_157;
      end
    end else begin
      buffer_4_pht_index <= _GEN_157;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_4_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h4 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_4_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_4_addr_misaligned <= _GEN_165;
      end
    end else begin
      buffer_4_addr_misaligned <= _GEN_165;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_4_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h4 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_4_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_4_access_fault <= _GEN_173;
      end
    end else begin
      buffer_4_access_fault <= _GEN_173;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_4_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h4 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_4_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_4_page_fault <= _GEN_181;
      end
    end else begin
      buffer_4_page_fault <= _GEN_181;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_4_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h4 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_4_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_4_pc <= _GEN_189;
      end
    end else begin
      buffer_4_pc <= _GEN_189;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_5_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h5 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_5_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_5_inst <= _GEN_150;
      end
    end else begin
      buffer_5_inst <= _GEN_150;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_5_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h5 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_5_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_5_pht_index <= _GEN_158;
      end
    end else begin
      buffer_5_pht_index <= _GEN_158;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_5_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h5 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_5_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_5_addr_misaligned <= _GEN_166;
      end
    end else begin
      buffer_5_addr_misaligned <= _GEN_166;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_5_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h5 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_5_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_5_access_fault <= _GEN_174;
      end
    end else begin
      buffer_5_access_fault <= _GEN_174;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_5_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h5 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_5_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_5_page_fault <= _GEN_182;
      end
    end else begin
      buffer_5_page_fault <= _GEN_182;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_5_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h5 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_5_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_5_pc <= _GEN_190;
      end
    end else begin
      buffer_5_pc <= _GEN_190;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_6_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h6 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_6_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_6_inst <= _GEN_151;
      end
    end else begin
      buffer_6_inst <= _GEN_151;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_6_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h6 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_6_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_6_pht_index <= _GEN_159;
      end
    end else begin
      buffer_6_pht_index <= _GEN_159;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_6_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h6 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_6_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_6_addr_misaligned <= _GEN_167;
      end
    end else begin
      buffer_6_addr_misaligned <= _GEN_167;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_6_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h6 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_6_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_6_access_fault <= _GEN_175;
      end
    end else begin
      buffer_6_access_fault <= _GEN_175;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_6_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h6 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_6_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_6_page_fault <= _GEN_183;
      end
    end else begin
      buffer_6_page_fault <= _GEN_183;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_6_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h6 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_6_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_6_pc <= _GEN_191;
      end
    end else begin
      buffer_6_pc <= _GEN_191;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_7_inst <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h7 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_7_inst <= io_write_1_inst; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_7_inst <= _GEN_152;
      end
    end else begin
      buffer_7_inst <= _GEN_152;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_7_pht_index <= 6'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h7 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_7_pht_index <= io_write_1_pht_index; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_7_pht_index <= _GEN_160;
      end
    end else begin
      buffer_7_pht_index <= _GEN_160;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_7_addr_misaligned <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h7 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_7_addr_misaligned <= io_write_1_addr_misaligned; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_7_addr_misaligned <= _GEN_168;
      end
    end else begin
      buffer_7_addr_misaligned <= _GEN_168;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_7_access_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h7 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_7_access_fault <= io_write_1_access_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_7_access_fault <= _GEN_176;
      end
    end else begin
      buffer_7_access_fault <= _GEN_176;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_7_page_fault <= 1'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h7 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_7_page_fault <= io_write_1_page_fault; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_7_page_fault <= _GEN_184;
      end
    end else begin
      buffer_7_page_fault <= _GEN_184;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
      buffer_7_pc <= 64'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 30:23]
    end else if (io_wen_1) begin // @[playground/src/pipeline/fetch/InstFifo.scala 83:21]
      if (3'h7 == _T_3) begin // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
        buffer_7_pc <= io_write_1_pc; // @[playground/src/pipeline/fetch/InstFifo.scala 84:29]
      end else begin
        buffer_7_pc <= _GEN_192;
      end
    end else begin
      buffer_7_pc <= _GEN_192;
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 33:24]
      enq_ptr <= 3'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 33:24]
    end else if (io_do_flush) begin // @[playground/src/pipeline/fetch/InstFifo.scala 88:21]
      enq_ptr <= 3'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 89:13]
    end else begin
      enq_ptr <= _enq_ptr_T_1; // @[playground/src/pipeline/fetch/InstFifo.scala 91:13]
    end
    if (reset) begin // @[playground/src/pipeline/fetch/InstFifo.scala 34:24]
      deq_ptr <= 3'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 34:24]
    end else if (io_do_flush) begin // @[playground/src/pipeline/fetch/InstFifo.scala 73:21]
      deq_ptr <= 3'h0; // @[playground/src/pipeline/fetch/InstFifo.scala 74:13]
    end else begin
      deq_ptr <= _deq_ptr_T_1; // @[playground/src/pipeline/fetch/InstFifo.scala 76:13]
    end
    count <= _GEN_297[2:0]; // @[playground/src/pipeline/fetch/InstFifo.scala 35:{24,24} 101:9]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  buffer_0_inst = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0_pht_index = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_0_addr_misaligned = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_0_access_fault = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_0_page_fault = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  buffer_0_pc = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  buffer_1_inst = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_1_pht_index = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_1_addr_misaligned = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_1_access_fault = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_1_page_fault = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  buffer_1_pc = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  buffer_2_inst = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_2_pht_index = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_2_addr_misaligned = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_2_access_fault = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_2_page_fault = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  buffer_2_pc = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  buffer_3_inst = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_3_pht_index = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_3_addr_misaligned = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_3_access_fault = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_3_page_fault = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  buffer_3_pc = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  buffer_4_inst = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_4_pht_index = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_4_addr_misaligned = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_4_access_fault = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_4_page_fault = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  buffer_4_pc = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  buffer_5_inst = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_5_pht_index = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_5_addr_misaligned = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_5_access_fault = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_5_page_fault = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  buffer_5_pc = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  buffer_6_inst = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_6_pht_index = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_6_addr_misaligned = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  buffer_6_access_fault = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_6_page_fault = _RAND_40[0:0];
  _RAND_41 = {2{`RANDOM}};
  buffer_6_pc = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  buffer_7_inst = _RAND_42[63:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_7_pht_index = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_7_addr_misaligned = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_7_access_fault = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_7_page_fault = _RAND_46[0:0];
  _RAND_47 = {2{`RANDOM}};
  buffer_7_pc = _RAND_47[63:0];
  _RAND_48 = {1{`RANDOM}};
  enq_ptr = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  deq_ptr = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  count = _RAND_50[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder(
  input  [63:0] io_in_inst, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output        io_out_info_inst_legal, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output        io_out_info_src1_ren, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [4:0]  io_out_info_src1_raddr, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output        io_out_info_src2_ren, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [4:0]  io_out_info_src2_raddr, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [2:0]  io_out_info_fusel, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [6:0]  io_out_info_op, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output        io_out_info_reg_wen, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [4:0]  io_out_info_reg_waddr, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [63:0] io_out_info_imm, // @[playground/src/pipeline/decode/Decoder.scala 9:14]
  output [63:0] io_out_info_inst // @[playground/src/pipeline/decode/Decoder.scala 9:14]
);
  wire [63:0] _T = io_in_inst & 64'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_1 = 64'h13 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_2 = io_in_inst & 64'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_3 = 64'h1013 == _T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_5 = 64'h2013 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_7 = 64'h3013 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_9 = 64'h4013 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_11 = 64'h5013 == _T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_13 = 64'h6013 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_15 = 64'h7013 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_17 = 64'h40005013 == _T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_18 = io_in_inst & 64'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_19 = 64'h33 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_21 = 64'h1033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_23 = 64'h2033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_25 = 64'h3033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_27 = 64'h4033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_29 = 64'h5033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_31 = 64'h6033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_33 = 64'h7033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_35 = 64'h40000033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_37 = 64'h40005033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_38 = io_in_inst & 64'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_39 = 64'h17 == _T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_41 = 64'h37 == _T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_43 = 64'h6f == _T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_45 = 64'h67 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_47 = 64'h63 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_49 = 64'h1063 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_51 = 64'h4063 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_53 = 64'h5063 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_55 = 64'h6063 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_57 = 64'h7063 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_59 = 64'h3 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_61 = 64'h1003 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_63 = 64'h2003 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_65 = 64'h4003 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_67 = 64'h5003 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_69 = 64'h23 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_71 = 64'h1023 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_73 = 64'h2023 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_75 = 64'h1b == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_77 = 64'h101b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_79 = 64'h501b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_81 = 64'h4000501b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_83 = 64'h103b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_85 = 64'h503b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_87 = 64'h4000503b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_89 = 64'h3b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_91 = 64'h4000003b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_93 = 64'h6003 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_95 = 64'h3003 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_97 = 64'h3023 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_99 = 64'h2000033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_101 = 64'h2001033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_103 = 64'h2002033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_105 = 64'h2003033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_107 = 64'h2004033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_109 = 64'h2005033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_111 = 64'h2006033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_113 = 64'h2007033 == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_115 = 64'h200003b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_117 = 64'h200403b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_119 = 64'h200503b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_121 = 64'h200603b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_123 = 64'h200703b == _T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_124 = io_in_inst & 64'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_125 = 64'h1000302f == _T_124; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_127 = 64'h1000202f == _T_124; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_128 = io_in_inst & 64'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_129 = 64'h1800302f == _T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_131 = 64'h1800202f == _T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_132 = io_in_inst & 64'hf800607f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_133 = 64'h800202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_135 = 64'h202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_137 = 64'h2000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_139 = 64'h6000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_141 = 64'h4000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_143 = 64'h8000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_145 = 64'ha000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_147 = 64'hc000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_149 = 64'he000202f == _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_150 = io_in_inst & 64'hffffffff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_151 = 64'h73 == _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_153 = 64'h100073 == _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_155 = 64'h30200073 == _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_157 = 64'hf == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_159 = 64'h10500073 == _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_161 = 64'h10200073 == _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _T_162 = io_in_inst & 64'hfe007fff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_163 = 64'h12000073 == _T_162; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_165 = 64'h1073 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_167 = 64'h2073 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_169 = 64'h3073 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_171 = 64'h5073 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_173 = 64'h6073 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_175 = 64'h7073 == _T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _T_177 = 64'h100f == _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _T_179 = _T_175 ? 3'h4 : {{2'd0}, _T_177}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_180 = _T_173 ? 3'h4 : _T_179; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_181 = _T_171 ? 3'h4 : _T_180; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_182 = _T_169 ? 3'h4 : _T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_183 = _T_167 ? 3'h4 : _T_182; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_184 = _T_165 ? 3'h4 : _T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_185 = _T_163 ? 3'h5 : _T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_186 = _T_161 ? 3'h4 : _T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_187 = _T_159 ? 3'h4 : _T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_188 = _T_157 ? 3'h2 : _T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_189 = _T_155 ? 3'h4 : _T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_190 = _T_153 ? 3'h4 : _T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_191 = _T_151 ? 3'h4 : _T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_192 = _T_149 ? 3'h5 : _T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_193 = _T_147 ? 3'h5 : _T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_194 = _T_145 ? 3'h5 : _T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_195 = _T_143 ? 3'h5 : _T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_196 = _T_141 ? 3'h5 : _T_195; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_197 = _T_139 ? 3'h5 : _T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_198 = _T_137 ? 3'h5 : _T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_199 = _T_135 ? 3'h5 : _T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_200 = _T_133 ? 3'h5 : _T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_201 = _T_131 ? 4'hf : {{1'd0}, _T_200}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_202 = _T_129 ? 4'hf : _T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_203 = _T_127 ? 4'h4 : _T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_204 = _T_125 ? 4'h4 : _T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_205 = _T_123 ? 4'h5 : _T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_206 = _T_121 ? 4'h5 : _T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_207 = _T_119 ? 4'h5 : _T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_208 = _T_117 ? 4'h5 : _T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_209 = _T_115 ? 4'h5 : _T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_210 = _T_113 ? 4'h5 : _T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_211 = _T_111 ? 4'h5 : _T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_212 = _T_109 ? 4'h5 : _T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_213 = _T_107 ? 4'h5 : _T_212; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_214 = _T_105 ? 4'h5 : _T_213; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_215 = _T_103 ? 4'h5 : _T_214; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_216 = _T_101 ? 4'h5 : _T_215; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_217 = _T_99 ? 4'h5 : _T_216; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_218 = _T_97 ? 4'h2 : _T_217; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_219 = _T_95 ? 4'h4 : _T_218; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_220 = _T_93 ? 4'h4 : _T_219; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_221 = _T_91 ? 4'h5 : _T_220; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_222 = _T_89 ? 4'h5 : _T_221; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_223 = _T_87 ? 4'h5 : _T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_224 = _T_85 ? 4'h5 : _T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_225 = _T_83 ? 4'h5 : _T_224; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_226 = _T_81 ? 4'h4 : _T_225; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_227 = _T_79 ? 4'h4 : _T_226; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_228 = _T_77 ? 4'h4 : _T_227; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_229 = _T_75 ? 4'h4 : _T_228; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_230 = _T_73 ? 4'h2 : _T_229; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_231 = _T_71 ? 4'h2 : _T_230; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_232 = _T_69 ? 4'h2 : _T_231; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_233 = _T_67 ? 4'h4 : _T_232; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_234 = _T_65 ? 4'h4 : _T_233; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_235 = _T_63 ? 4'h4 : _T_234; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_236 = _T_61 ? 4'h4 : _T_235; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_237 = _T_59 ? 4'h4 : _T_236; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_238 = _T_57 ? 4'h1 : _T_237; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_239 = _T_55 ? 4'h1 : _T_238; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_240 = _T_53 ? 4'h1 : _T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_241 = _T_51 ? 4'h1 : _T_240; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_242 = _T_49 ? 4'h1 : _T_241; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_243 = _T_47 ? 4'h1 : _T_242; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_244 = _T_45 ? 4'h4 : _T_243; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_245 = _T_43 ? 4'h7 : _T_244; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_246 = _T_41 ? 4'h6 : _T_245; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_247 = _T_39 ? 4'h6 : _T_246; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_248 = _T_37 ? 4'h5 : _T_247; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_249 = _T_35 ? 4'h5 : _T_248; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_250 = _T_33 ? 4'h5 : _T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_251 = _T_31 ? 4'h5 : _T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_252 = _T_29 ? 4'h5 : _T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_253 = _T_27 ? 4'h5 : _T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_254 = _T_25 ? 4'h5 : _T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_255 = _T_23 ? 4'h5 : _T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_256 = _T_21 ? 4'h5 : _T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_257 = _T_19 ? 4'h5 : _T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_258 = _T_17 ? 4'h4 : _T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_259 = _T_15 ? 4'h4 : _T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_260 = _T_13 ? 4'h4 : _T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_261 = _T_11 ? 4'h4 : _T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_262 = _T_9 ? 4'h4 : _T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_263 = _T_7 ? 4'h4 : _T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_264 = _T_5 ? 4'h4 : _T_263; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_265 = _T_3 ? 4'h4 : _T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] instrType = _T_1 ? 4'h4 : _T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_266 = _T_177 ? 3'h4 : 3'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_267 = _T_175 ? 3'h3 : _T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_268 = _T_173 ? 3'h3 : _T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_269 = _T_171 ? 3'h3 : _T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_270 = _T_169 ? 3'h3 : _T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_271 = _T_167 ? 3'h3 : _T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_272 = _T_165 ? 3'h3 : _T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_273 = _T_163 ? 3'h4 : _T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_274 = _T_161 ? 3'h3 : _T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_275 = _T_159 ? 3'h0 : _T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_276 = _T_157 ? 3'h4 : _T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_277 = _T_155 ? 3'h3 : _T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_278 = _T_153 ? 3'h3 : _T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_279 = _T_151 ? 3'h3 : _T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_280 = _T_149 ? 3'h1 : _T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_281 = _T_147 ? 3'h1 : _T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_282 = _T_145 ? 3'h1 : _T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_283 = _T_143 ? 3'h1 : _T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_284 = _T_141 ? 3'h1 : _T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_285 = _T_139 ? 3'h1 : _T_284; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_286 = _T_137 ? 3'h1 : _T_285; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_287 = _T_135 ? 3'h1 : _T_286; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_288 = _T_133 ? 3'h1 : _T_287; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_289 = _T_131 ? 3'h1 : _T_288; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_290 = _T_129 ? 3'h1 : _T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_291 = _T_127 ? 3'h1 : _T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_292 = _T_125 ? 3'h1 : _T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_293 = _T_123 ? 3'h2 : _T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_294 = _T_121 ? 3'h2 : _T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_295 = _T_119 ? 3'h2 : _T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_296 = _T_117 ? 3'h2 : _T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_297 = _T_115 ? 3'h2 : _T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_298 = _T_113 ? 3'h2 : _T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_299 = _T_111 ? 3'h2 : _T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_300 = _T_109 ? 3'h2 : _T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_301 = _T_107 ? 3'h2 : _T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_302 = _T_105 ? 3'h2 : _T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_303 = _T_103 ? 3'h2 : _T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_304 = _T_101 ? 3'h2 : _T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_305 = _T_99 ? 3'h2 : _T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_306 = _T_97 ? 3'h1 : _T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_307 = _T_95 ? 3'h1 : _T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_308 = _T_93 ? 3'h1 : _T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_309 = _T_91 ? 3'h0 : _T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_310 = _T_89 ? 3'h0 : _T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_311 = _T_87 ? 3'h0 : _T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_312 = _T_85 ? 3'h0 : _T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_313 = _T_83 ? 3'h0 : _T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_314 = _T_81 ? 3'h0 : _T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_315 = _T_79 ? 3'h0 : _T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_316 = _T_77 ? 3'h0 : _T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_317 = _T_75 ? 3'h0 : _T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_318 = _T_73 ? 3'h1 : _T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_319 = _T_71 ? 3'h1 : _T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_320 = _T_69 ? 3'h1 : _T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_321 = _T_67 ? 3'h1 : _T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_322 = _T_65 ? 3'h1 : _T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_323 = _T_63 ? 3'h1 : _T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_324 = _T_61 ? 3'h1 : _T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_325 = _T_59 ? 3'h1 : _T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_326 = _T_57 ? 3'h5 : _T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_327 = _T_55 ? 3'h5 : _T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_328 = _T_53 ? 3'h5 : _T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_329 = _T_51 ? 3'h5 : _T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_330 = _T_49 ? 3'h5 : _T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_331 = _T_47 ? 3'h5 : _T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_332 = _T_45 ? 3'h5 : _T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_333 = _T_43 ? 3'h5 : _T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_334 = _T_41 ? 3'h0 : _T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_335 = _T_39 ? 3'h0 : _T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_336 = _T_37 ? 3'h0 : _T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_337 = _T_35 ? 3'h0 : _T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_338 = _T_33 ? 3'h0 : _T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_339 = _T_31 ? 3'h0 : _T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_340 = _T_29 ? 3'h0 : _T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_341 = _T_27 ? 3'h0 : _T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_342 = _T_25 ? 3'h0 : _T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_343 = _T_23 ? 3'h0 : _T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_344 = _T_21 ? 3'h0 : _T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_345 = _T_19 ? 3'h0 : _T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_346 = _T_17 ? 3'h0 : _T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_347 = _T_15 ? 3'h0 : _T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_348 = _T_13 ? 3'h0 : _T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_349 = _T_11 ? 3'h0 : _T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_350 = _T_9 ? 3'h0 : _T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_351 = _T_7 ? 3'h0 : _T_350; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_352 = _T_5 ? 3'h0 : _T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_353 = _T_3 ? 3'h0 : _T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_354 = _T_177 ? 6'h1 : 6'h20; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_355 = _T_175 ? 6'h7 : _T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_356 = _T_173 ? 6'h6 : _T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_357 = _T_171 ? 6'h5 : _T_356; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_358 = _T_169 ? 6'h3 : _T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_359 = _T_167 ? 6'h2 : _T_358; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_360 = _T_165 ? 6'h1 : _T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_361 = _T_163 ? 6'h2 : _T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_362 = _T_161 ? 6'hb : _T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_363 = _T_159 ? 6'h20 : _T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_364 = _T_157 ? 6'h0 : _T_363; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_365 = _T_155 ? 6'ha : _T_364; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_366 = _T_153 ? 6'h9 : _T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_367 = _T_151 ? 6'h8 : _T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_368 = _T_149 ? 6'h32 : _T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_369 = _T_147 ? 6'h31 : _T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_370 = _T_145 ? 6'h30 : _T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_371 = _T_143 ? 6'h37 : _T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_372 = _T_141 ? 6'h26 : _T_371; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_373 = _T_139 ? 6'h25 : _T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _T_374 = _T_137 ? 6'h24 : _T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_375 = _T_135 ? 7'h63 : {{1'd0}, _T_374}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_376 = _T_133 ? 7'h22 : _T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_377 = _T_131 ? 7'h21 : _T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_378 = _T_129 ? 7'h21 : _T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_379 = _T_127 ? 7'h20 : _T_378; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_380 = _T_125 ? 7'h20 : _T_379; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_381 = _T_123 ? 7'hf : _T_380; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_382 = _T_121 ? 7'he : _T_381; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_383 = _T_119 ? 7'hd : _T_382; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_384 = _T_117 ? 7'hc : _T_383; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_385 = _T_115 ? 7'h8 : _T_384; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_386 = _T_113 ? 7'h7 : _T_385; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_387 = _T_111 ? 7'h6 : _T_386; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_388 = _T_109 ? 7'h5 : _T_387; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_389 = _T_107 ? 7'h4 : _T_388; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_390 = _T_105 ? 7'h3 : _T_389; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_391 = _T_103 ? 7'h2 : _T_390; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_392 = _T_101 ? 7'h1 : _T_391; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_393 = _T_99 ? 7'h0 : _T_392; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_394 = _T_97 ? 7'hb : _T_393; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_395 = _T_95 ? 7'h3 : _T_394; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_396 = _T_93 ? 7'h6 : _T_395; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_397 = _T_91 ? 7'h18 : _T_396; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_398 = _T_89 ? 7'h30 : _T_397; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_399 = _T_87 ? 7'h1d : _T_398; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_400 = _T_85 ? 7'h15 : _T_399; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_401 = _T_83 ? 7'h11 : _T_400; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_402 = _T_81 ? 7'h1d : _T_401; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_403 = _T_79 ? 7'h15 : _T_402; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_404 = _T_77 ? 7'h11 : _T_403; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_405 = _T_75 ? 7'h30 : _T_404; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_406 = _T_73 ? 7'ha : _T_405; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_407 = _T_71 ? 7'h9 : _T_406; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_408 = _T_69 ? 7'h8 : _T_407; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_409 = _T_67 ? 7'h5 : _T_408; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_410 = _T_65 ? 7'h4 : _T_409; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_411 = _T_63 ? 7'h2 : _T_410; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_412 = _T_61 ? 7'h1 : _T_411; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_413 = _T_59 ? 7'h0 : _T_412; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_414 = _T_57 ? 7'h7 : _T_413; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_415 = _T_55 ? 7'h6 : _T_414; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_416 = _T_53 ? 7'h5 : _T_415; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_417 = _T_51 ? 7'h4 : _T_416; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_418 = _T_49 ? 7'h1 : _T_417; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_419 = _T_47 ? 7'h0 : _T_418; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_420 = _T_45 ? 7'ha : _T_419; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_421 = _T_43 ? 7'h8 : _T_420; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_422 = _T_41 ? 7'h20 : _T_421; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_423 = _T_39 ? 7'h20 : _T_422; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_424 = _T_37 ? 7'hd : _T_423; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_425 = _T_35 ? 7'h8 : _T_424; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_426 = _T_33 ? 7'h7 : _T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_427 = _T_31 ? 7'h6 : _T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_428 = _T_29 ? 7'h5 : _T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_429 = _T_27 ? 7'h4 : _T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_430 = _T_25 ? 7'h3 : _T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_431 = _T_23 ? 7'h2 : _T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_432 = _T_21 ? 7'h1 : _T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_433 = _T_19 ? 7'h20 : _T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_434 = _T_17 ? 7'hd : _T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_435 = _T_15 ? 7'h7 : _T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_436 = _T_13 ? 7'h6 : _T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_437 = _T_11 ? 7'h5 : _T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_438 = _T_9 ? 7'h4 : _T_437; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_439 = _T_7 ? 7'h3 : _T_438; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_440 = _T_5 ? 7'h2 : _T_439; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _T_441 = _T_3 ? 7'h1 : _T_440; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _src1Type_T = 4'h4 == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  _src1Type_T_2 = 4'h2 == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  _src1Type_T_3 = 4'hf == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  _src1Type_T_4 = 4'h1 == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  _src1Type_T_5 = 4'h6 == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  _src1Type_T_6 = 4'h7 == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  _src1Type_T_7 = 4'h0 == instrType; // @[playground/src/defines/Util.scala 46:34]
  wire  src1Type = _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rs = io_in_inst[19:15]; // @[playground/src/pipeline/decode/Decoder.scala 37:27]
  wire [4:0] rt = io_in_inst[24:20]; // @[playground/src/pipeline/decode/Decoder.scala 37:41]
  wire [4:0] rd = io_in_inst[11:7]; // @[playground/src/pipeline/decode/Decoder.scala 37:55]
  wire  io_out_info_imm_signBit = io_in_inst[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [51:0] _io_out_info_imm_T_2 = io_out_info_imm_signBit ? 52'hfffffffffffff : 52'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_out_info_imm_T_3 = {_io_out_info_imm_T_2,io_in_inst[31:20]}; // @[playground/src/defines/Util.scala 34:44]
  wire [11:0] _io_out_info_imm_T_6 = {io_in_inst[31:25],rd}; // @[playground/src/pipeline/decode/Decoder.scala 54:34]
  wire  io_out_info_imm_signBit_1 = _io_out_info_imm_T_6[11]; // @[playground/src/defines/Util.scala 33:20]
  wire [51:0] _io_out_info_imm_T_8 = io_out_info_imm_signBit_1 ? 52'hfffffffffffff : 52'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_out_info_imm_T_9 = {_io_out_info_imm_T_8,io_in_inst[31:25],rd}; // @[playground/src/defines/Util.scala 34:44]
  wire [12:0] _io_out_info_imm_T_20 = {io_in_inst[31],io_in_inst[7],io_in_inst[30:25],io_in_inst[11:8],1'h0}; // @[playground/src/pipeline/decode/Decoder.scala 56:34]
  wire  io_out_info_imm_signBit_3 = _io_out_info_imm_T_20[12]; // @[playground/src/defines/Util.scala 33:20]
  wire [50:0] _io_out_info_imm_T_22 = io_out_info_imm_signBit_3 ? 51'h7ffffffffffff : 51'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_out_info_imm_T_23 = {_io_out_info_imm_T_22,io_in_inst[31],io_in_inst[7],io_in_inst[30:25],io_in_inst[
    11:8],1'h0}; // @[playground/src/defines/Util.scala 34:44]
  wire [31:0] _io_out_info_imm_T_25 = {io_in_inst[31:12],12'h0}; // @[playground/src/pipeline/decode/Decoder.scala 57:34]
  wire  io_out_info_imm_signBit_4 = _io_out_info_imm_T_25[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _io_out_info_imm_T_27 = io_out_info_imm_signBit_4 ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_out_info_imm_T_28 = {_io_out_info_imm_T_27,io_in_inst[31:12],12'h0}; // @[playground/src/defines/Util.scala 34:44]
  wire [20:0] _io_out_info_imm_T_33 = {io_in_inst[31],io_in_inst[19:12],io_in_inst[20],io_in_inst[30:21],1'h0}; // @[playground/src/pipeline/decode/Decoder.scala 58:34]
  wire  io_out_info_imm_signBit_5 = _io_out_info_imm_T_33[20]; // @[playground/src/defines/Util.scala 33:20]
  wire [42:0] _io_out_info_imm_T_35 = io_out_info_imm_signBit_5 ? 43'h7ffffffffff : 43'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_out_info_imm_T_36 = {_io_out_info_imm_T_35,io_in_inst[31],io_in_inst[19:12],io_in_inst[20],io_in_inst[
    30:21],1'h0}; // @[playground/src/defines/Util.scala 34:44]
  wire [63:0] _io_out_info_imm_T_43 = _src1Type_T ? _io_out_info_imm_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_44 = _src1Type_T_2 ? _io_out_info_imm_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_45 = _src1Type_T_3 ? _io_out_info_imm_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_46 = _src1Type_T_4 ? _io_out_info_imm_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_47 = _src1Type_T_5 ? _io_out_info_imm_T_28 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_48 = _src1Type_T_6 ? _io_out_info_imm_T_36 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_49 = _io_out_info_imm_T_43 | _io_out_info_imm_T_44; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_50 = _io_out_info_imm_T_49 | _io_out_info_imm_T_45; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_51 = _io_out_info_imm_T_50 | _io_out_info_imm_T_46; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_info_imm_T_52 = _io_out_info_imm_T_51 | _io_out_info_imm_T_47; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_info_inst_legal = instrType != 4'h0; // @[playground/src/pipeline/decode/Decoder.scala 41:39]
  assign io_out_info_src1_ren = ~src1Type; // @[playground/src/pipeline/decode/Decoder.scala 42:38]
  assign io_out_info_src1_raddr = io_out_info_src1_ren ? rs : 5'h0; // @[playground/src/pipeline/decode/Decoder.scala 43:32]
  assign io_out_info_src2_ren = ~src2Type; // @[playground/src/pipeline/decode/Decoder.scala 44:38]
  assign io_out_info_src2_raddr = io_out_info_src2_ren ? rt : 5'h0; // @[playground/src/pipeline/decode/Decoder.scala 45:32]
  assign io_out_info_fusel = _T_1 ? 3'h0 : _T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  assign io_out_info_op = _T_1 ? 7'h20 : _T_441; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  assign io_out_info_reg_wen = instrType[2]; // @[playground/src/defines/isa/Instructions.scala 16:50]
  assign io_out_info_reg_waddr = instrType[2] ? rd : 5'h0; // @[playground/src/pipeline/decode/Decoder.scala 49:32]
  assign io_out_info_imm = _io_out_info_imm_T_52 | _io_out_info_imm_T_48; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_info_inst = io_in_inst; // @[playground/src/pipeline/decode/Decoder.scala 40:26]
endmodule
module JumpCtrl(
  input         io_in_info_valid, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [4:0]  io_in_info_src1_raddr, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [2:0]  io_in_info_fusel, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [6:0]  io_in_info_op, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [63:0] io_in_src_info_src1_data, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [63:0] io_in_src_info_src2_data, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input         io_in_forward_0_exe_wen, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [4:0]  io_in_forward_0_exe_waddr, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input         io_in_forward_0_mem_wen, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [4:0]  io_in_forward_0_mem_waddr, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input         io_in_forward_1_exe_wen, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [4:0]  io_in_forward_1_exe_waddr, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input         io_in_forward_1_mem_wen, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  input  [4:0]  io_in_forward_1_mem_waddr, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  output        io_out_jump_register, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  output        io_out_jump, // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
  output [63:0] io_out_jump_target // @[playground/src/pipeline/decode/JumpCtrl.scala 11:14]
);
  wire  _jump_inst_T_2 = io_in_info_fusel == 3'h5; // @[playground/src/pipeline/decode/JumpCtrl.scala 28:73]
  wire  jump_inst = 7'h8 == io_in_info_op & io_in_info_fusel == 3'h5; // @[playground/src/pipeline/decode/JumpCtrl.scala 28:64]
  wire  jump_register_inst = 7'ha == io_in_info_op & _jump_inst_T_2; // @[playground/src/pipeline/decode/JumpCtrl.scala 29:65]
  wire  _io_out_jump_register_T_5 = io_in_forward_1_exe_wen & io_in_info_src1_raddr == io_in_forward_1_exe_waddr; // @[playground/src/pipeline/decode/JumpCtrl.scala 34:31]
  wire  _io_out_jump_register_T_6 = io_in_forward_0_exe_wen & io_in_info_src1_raddr == io_in_forward_0_exe_waddr |
    _io_out_jump_register_T_5; // @[playground/src/pipeline/decode/JumpCtrl.scala 33:89]
  wire  _io_out_jump_register_T_8 = io_in_forward_0_mem_wen & io_in_info_src1_raddr == io_in_forward_0_mem_waddr; // @[playground/src/pipeline/decode/JumpCtrl.scala 35:31]
  wire  _io_out_jump_register_T_9 = _io_out_jump_register_T_6 | _io_out_jump_register_T_8; // @[playground/src/pipeline/decode/JumpCtrl.scala 34:88]
  wire  _io_out_jump_register_T_11 = io_in_forward_1_mem_wen & io_in_info_src1_raddr == io_in_forward_1_mem_waddr; // @[playground/src/pipeline/decode/JumpCtrl.scala 36:31]
  wire  _io_out_jump_register_T_12 = _io_out_jump_register_T_9 | _io_out_jump_register_T_11; // @[playground/src/pipeline/decode/JumpCtrl.scala 35:88]
  wire [63:0] _io_out_jump_target_T_1 = io_in_src_info_src1_data + io_in_src_info_src2_data; // @[playground/src/pipeline/decode/JumpCtrl.scala 45:30]
  wire [63:0] _io_out_jump_target_T_5 = _io_out_jump_target_T_1 & 64'hfffffffffffffffe; // @[playground/src/pipeline/decode/JumpCtrl.scala 46:59]
  assign io_out_jump_register = jump_register_inst & |io_in_info_src1_raddr & _io_out_jump_register_T_12; // @[playground/src/pipeline/decode/JumpCtrl.scala 32:77]
  assign io_out_jump = (jump_inst | jump_register_inst & ~io_out_jump_register) & io_in_info_valid; // @[playground/src/pipeline/decode/JumpCtrl.scala 30:77]
  assign io_out_jump_target = jump_inst ? _io_out_jump_target_T_1 : _io_out_jump_target_T_5; // @[playground/src/pipeline/decode/JumpCtrl.scala 43:28]
endmodule
module ForwardCtrl(
  input         io_in_forward_0_exe_wen, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_forward_0_exe_waddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_forward_0_exe_wdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input         io_in_forward_0_is_load, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input         io_in_forward_0_mem_wen, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_forward_0_mem_waddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_forward_0_mem_wdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input         io_in_forward_1_exe_wen, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_forward_1_exe_waddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_forward_1_exe_wdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input         io_in_forward_1_is_load, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input         io_in_forward_1_mem_wen, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_forward_1_mem_waddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_forward_1_mem_wdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_regfile_0_src1_raddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_regfile_0_src1_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_regfile_0_src2_raddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_regfile_0_src2_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_regfile_1_src1_raddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_regfile_1_src1_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [4:0]  io_in_regfile_1_src2_raddr, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  input  [63:0] io_in_regfile_1_src2_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  output [63:0] io_out_inst_0_src1_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  output [63:0] io_out_inst_0_src2_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  output [63:0] io_out_inst_1_src1_rdata, // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
  output [63:0] io_out_inst_1_src2_rdata // @[playground/src/pipeline/decode/ForwardCtrl.scala 11:14]
);
  wire  _T = io_in_forward_0_mem_waddr == io_in_regfile_0_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 34:38]
  wire  _T_1 = io_in_forward_0_mem_wen & _T; // @[playground/src/pipeline/decode/ForwardCtrl.scala 33:34]
  wire [63:0] _GEN_0 = _T_1 ? io_in_forward_0_mem_wdata : io_in_regfile_0_src1_rdata; // @[playground/src/pipeline/decode/ForwardCtrl.scala 25:31 35:9 36:35]
  wire  _T_2 = io_in_forward_0_mem_waddr == io_in_regfile_0_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 40:38]
  wire  _T_3 = io_in_forward_0_mem_wen & _T_2; // @[playground/src/pipeline/decode/ForwardCtrl.scala 39:34]
  wire [63:0] _GEN_1 = _T_3 ? io_in_forward_0_mem_wdata : io_in_regfile_0_src2_rdata; // @[playground/src/pipeline/decode/ForwardCtrl.scala 26:31 41:9 42:35]
  wire  _T_4 = io_in_forward_1_mem_waddr == io_in_regfile_0_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 34:38]
  wire  _T_5 = io_in_forward_1_mem_wen & _T_4; // @[playground/src/pipeline/decode/ForwardCtrl.scala 33:34]
  wire [63:0] _GEN_2 = _T_5 ? io_in_forward_1_mem_wdata : _GEN_0; // @[playground/src/pipeline/decode/ForwardCtrl.scala 35:9 36:35]
  wire  _T_6 = io_in_forward_1_mem_waddr == io_in_regfile_0_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 40:38]
  wire  _T_7 = io_in_forward_1_mem_wen & _T_6; // @[playground/src/pipeline/decode/ForwardCtrl.scala 39:34]
  wire [63:0] _GEN_3 = _T_7 ? io_in_forward_1_mem_wdata : _GEN_1; // @[playground/src/pipeline/decode/ForwardCtrl.scala 41:9 42:35]
  wire  _T_8 = io_in_forward_0_mem_waddr == io_in_regfile_1_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 34:38]
  wire  _T_9 = io_in_forward_0_mem_wen & _T_8; // @[playground/src/pipeline/decode/ForwardCtrl.scala 33:34]
  wire [63:0] _GEN_4 = _T_9 ? io_in_forward_0_mem_wdata : io_in_regfile_1_src1_rdata; // @[playground/src/pipeline/decode/ForwardCtrl.scala 25:31 35:9 36:35]
  wire  _T_10 = io_in_forward_0_mem_waddr == io_in_regfile_1_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 40:38]
  wire  _T_11 = io_in_forward_0_mem_wen & _T_10; // @[playground/src/pipeline/decode/ForwardCtrl.scala 39:34]
  wire [63:0] _GEN_5 = _T_11 ? io_in_forward_0_mem_wdata : io_in_regfile_1_src2_rdata; // @[playground/src/pipeline/decode/ForwardCtrl.scala 26:31 41:9 42:35]
  wire  _T_12 = io_in_forward_1_mem_waddr == io_in_regfile_1_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 34:38]
  wire  _T_13 = io_in_forward_1_mem_wen & _T_12; // @[playground/src/pipeline/decode/ForwardCtrl.scala 33:34]
  wire [63:0] _GEN_6 = _T_13 ? io_in_forward_1_mem_wdata : _GEN_4; // @[playground/src/pipeline/decode/ForwardCtrl.scala 35:9 36:35]
  wire  _T_14 = io_in_forward_1_mem_waddr == io_in_regfile_1_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 40:38]
  wire  _T_15 = io_in_forward_1_mem_wen & _T_14; // @[playground/src/pipeline/decode/ForwardCtrl.scala 39:34]
  wire [63:0] _GEN_7 = _T_15 ? io_in_forward_1_mem_wdata : _GEN_5; // @[playground/src/pipeline/decode/ForwardCtrl.scala 41:9 42:35]
  wire  _T_17 = io_in_forward_0_exe_wen & ~io_in_forward_0_is_load; // @[playground/src/pipeline/decode/ForwardCtrl.scala 51:34]
  wire  _T_18 = io_in_forward_0_exe_waddr == io_in_regfile_0_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 52:38]
  wire  _T_19 = io_in_forward_0_exe_wen & ~io_in_forward_0_is_load & _T_18; // @[playground/src/pipeline/decode/ForwardCtrl.scala 51:63]
  wire [63:0] _GEN_8 = _T_19 ? io_in_forward_0_exe_wdata : _GEN_2; // @[playground/src/pipeline/decode/ForwardCtrl.scala 53:9 54:35]
  wire  _T_22 = io_in_forward_0_exe_waddr == io_in_regfile_0_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 58:38]
  wire  _T_23 = _T_17 & _T_22; // @[playground/src/pipeline/decode/ForwardCtrl.scala 57:63]
  wire [63:0] _GEN_9 = _T_23 ? io_in_forward_0_exe_wdata : _GEN_3; // @[playground/src/pipeline/decode/ForwardCtrl.scala 59:9 60:35]
  wire  _T_25 = io_in_forward_1_exe_wen & ~io_in_forward_1_is_load; // @[playground/src/pipeline/decode/ForwardCtrl.scala 51:34]
  wire  _T_26 = io_in_forward_1_exe_waddr == io_in_regfile_0_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 52:38]
  wire  _T_27 = io_in_forward_1_exe_wen & ~io_in_forward_1_is_load & _T_26; // @[playground/src/pipeline/decode/ForwardCtrl.scala 51:63]
  wire [63:0] _GEN_10 = _T_27 ? io_in_forward_1_exe_wdata : _GEN_8; // @[playground/src/pipeline/decode/ForwardCtrl.scala 53:9 54:35]
  wire  _T_30 = io_in_forward_1_exe_waddr == io_in_regfile_0_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 58:38]
  wire  _T_31 = _T_25 & _T_30; // @[playground/src/pipeline/decode/ForwardCtrl.scala 57:63]
  wire [63:0] _GEN_11 = _T_31 ? io_in_forward_1_exe_wdata : _GEN_9; // @[playground/src/pipeline/decode/ForwardCtrl.scala 59:9 60:35]
  wire  _T_34 = io_in_forward_0_exe_waddr == io_in_regfile_1_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 52:38]
  wire  _T_35 = io_in_forward_0_exe_wen & ~io_in_forward_0_is_load & _T_34; // @[playground/src/pipeline/decode/ForwardCtrl.scala 51:63]
  wire [63:0] _GEN_12 = _T_35 ? io_in_forward_0_exe_wdata : _GEN_6; // @[playground/src/pipeline/decode/ForwardCtrl.scala 53:9 54:35]
  wire  _T_38 = io_in_forward_0_exe_waddr == io_in_regfile_1_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 58:38]
  wire  _T_39 = _T_17 & _T_38; // @[playground/src/pipeline/decode/ForwardCtrl.scala 57:63]
  wire [63:0] _GEN_13 = _T_39 ? io_in_forward_0_exe_wdata : _GEN_7; // @[playground/src/pipeline/decode/ForwardCtrl.scala 59:9 60:35]
  wire  _T_42 = io_in_forward_1_exe_waddr == io_in_regfile_1_src1_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 52:38]
  wire  _T_43 = io_in_forward_1_exe_wen & ~io_in_forward_1_is_load & _T_42; // @[playground/src/pipeline/decode/ForwardCtrl.scala 51:63]
  wire [63:0] _GEN_14 = _T_43 ? io_in_forward_1_exe_wdata : _GEN_12; // @[playground/src/pipeline/decode/ForwardCtrl.scala 53:9 54:35]
  wire  _T_46 = io_in_forward_1_exe_waddr == io_in_regfile_1_src2_raddr; // @[playground/src/pipeline/decode/ForwardCtrl.scala 58:38]
  wire  _T_47 = _T_25 & _T_46; // @[playground/src/pipeline/decode/ForwardCtrl.scala 57:63]
  wire [63:0] _GEN_15 = _T_47 ? io_in_forward_1_exe_wdata : _GEN_13; // @[playground/src/pipeline/decode/ForwardCtrl.scala 59:9 60:35]
  assign io_out_inst_0_src1_rdata = io_in_regfile_0_src1_raddr == 5'h0 ? 64'h0 : _GEN_10; // @[playground/src/pipeline/decode/ForwardCtrl.scala 67:47 68:33]
  assign io_out_inst_0_src2_rdata = io_in_regfile_0_src2_raddr == 5'h0 ? 64'h0 : _GEN_11; // @[playground/src/pipeline/decode/ForwardCtrl.scala 70:47 71:33]
  assign io_out_inst_1_src1_rdata = io_in_regfile_1_src1_raddr == 5'h0 ? 64'h0 : _GEN_14; // @[playground/src/pipeline/decode/ForwardCtrl.scala 67:47 68:33]
  assign io_out_inst_1_src2_rdata = io_in_regfile_1_src2_raddr == 5'h0 ? 64'h0 : _GEN_15; // @[playground/src/pipeline/decode/ForwardCtrl.scala 70:47 71:33]
endmodule
module Issue(
  input         io_allow_to_go, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_instFifo_empty, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_instFifo_almost_empty, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [2:0]  io_decodeInst_0_fusel, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [6:0]  io_decodeInst_0_op, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_decodeInst_0_reg_wen, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [4:0]  io_decodeInst_0_reg_waddr, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [63:0] io_decodeInst_0_inst, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_decodeInst_1_src1_ren, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [4:0]  io_decodeInst_1_src1_raddr, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_decodeInst_1_src2_ren, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [4:0]  io_decodeInst_1_src2_raddr, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [2:0]  io_decodeInst_1_fusel, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [6:0]  io_decodeInst_1_op, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [63:0] io_decodeInst_1_inst, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_execute_0_is_load, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [4:0]  io_execute_0_reg_waddr, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input         io_execute_1_is_load, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  input  [4:0]  io_execute_1_reg_waddr, // @[playground/src/pipeline/decode/Issue.scala 11:14]
  output        io_inst1_allow_to_go // @[playground/src/pipeline/decode/Issue.scala 11:14]
);
  wire  instFifo_invalid = io_instFifo_empty | io_instFifo_almost_empty; // @[playground/src/pipeline/decode/Issue.scala 30:46]
  wire  lsu_conflict = io_decodeInst_0_fusel == 3'h1 & io_decodeInst_1_fusel == 3'h1; // @[playground/src/pipeline/decode/Issue.scala 33:69]
  wire  mdu_conflict = io_decodeInst_0_fusel == 3'h2 & io_decodeInst_1_fusel == 3'h2; // @[playground/src/pipeline/decode/Issue.scala 34:69]
  wire  _csr_conflict_T = io_decodeInst_0_fusel == 3'h3; // @[playground/src/pipeline/decode/Issue.scala 35:44]
  wire  _csr_conflict_T_1 = io_decodeInst_1_fusel == 3'h3; // @[playground/src/pipeline/decode/Issue.scala 35:44]
  wire  csr_conflict = io_decodeInst_0_fusel == 3'h3 & io_decodeInst_1_fusel == 3'h3; // @[playground/src/pipeline/decode/Issue.scala 35:69]
  wire  struct_conflict = lsu_conflict | mdu_conflict | csr_conflict; // @[playground/src/pipeline/decode/Issue.scala 36:56]
  wire  _load_stall_T_5 = io_decodeInst_1_src2_ren & io_decodeInst_1_src2_raddr == io_execute_0_reg_waddr; // @[playground/src/pipeline/decode/Issue.scala 42:28]
  wire  _load_stall_T_6 = io_decodeInst_1_src1_ren & io_decodeInst_1_src1_raddr == io_execute_0_reg_waddr |
    _load_stall_T_5; // @[playground/src/pipeline/decode/Issue.scala 41:77]
  wire  _load_stall_T_7 = io_execute_0_is_load & |io_execute_0_reg_waddr & _load_stall_T_6; // @[playground/src/pipeline/decode/Issue.scala 40:60]
  wire  _load_stall_T_13 = io_decodeInst_1_src2_ren & io_decodeInst_1_src2_raddr == io_execute_1_reg_waddr; // @[playground/src/pipeline/decode/Issue.scala 45:30]
  wire  _load_stall_T_14 = io_decodeInst_1_src1_ren & io_decodeInst_1_src1_raddr == io_execute_1_reg_waddr |
    _load_stall_T_13; // @[playground/src/pipeline/decode/Issue.scala 44:79]
  wire  _load_stall_T_15 = io_execute_1_is_load & |io_execute_1_reg_waddr & _load_stall_T_14; // @[playground/src/pipeline/decode/Issue.scala 43:62]
  wire  load_stall = _load_stall_T_7 | _load_stall_T_15; // @[playground/src/pipeline/decode/Issue.scala 42:79]
  wire  _raw_reg_T_5 = io_decodeInst_0_reg_waddr == io_decodeInst_1_src2_raddr & io_decodeInst_1_src2_ren; // @[playground/src/pipeline/decode/Issue.scala 49:52]
  wire  _raw_reg_T_6 = io_decodeInst_0_reg_waddr == io_decodeInst_1_src1_raddr & io_decodeInst_1_src1_ren | _raw_reg_T_5
    ; // @[playground/src/pipeline/decode/Issue.scala 48:71]
  wire  raw_reg = io_decodeInst_0_reg_wen & |io_decodeInst_0_reg_waddr & _raw_reg_T_6; // @[playground/src/pipeline/decode/Issue.scala 47:48]
  wire  data_conflict = raw_reg | load_stall; // @[playground/src/pipeline/decode/Issue.scala 50:33]
  wire  is_bru = io_decodeInst_0_fusel == 3'h5 | io_decodeInst_1_fusel == 3'h5; // @[playground/src/pipeline/decode/Issue.scala 53:60]
  wire  is_mou = io_decodeInst_0_fusel == 3'h4 | io_decodeInst_1_fusel == 3'h4; // @[playground/src/pipeline/decode/Issue.scala 56:60]
  wire  _write_satp_T_2 = ~io_decodeInst_0_op[3]; // @[playground/src/defines/isa/Instructions.scala 159:27]
  wire  _write_satp_T_6 = _csr_conflict_T & _write_satp_T_2 & io_decodeInst_0_inst[31:20] == 12'h180; // @[playground/src/pipeline/decode/Issue.scala 61:71]
  wire  _write_satp_T_9 = ~io_decodeInst_1_op[3]; // @[playground/src/defines/isa/Instructions.scala 159:27]
  wire  _write_satp_T_13 = _csr_conflict_T_1 & _write_satp_T_9 & io_decodeInst_1_inst[31:20] == 12'h180; // @[playground/src/pipeline/decode/Issue.scala 61:71]
  wire [1:0] _write_satp_T_14 = {_write_satp_T_13,_write_satp_T_6}; // @[playground/src/pipeline/decode/Issue.scala 63:7]
  wire  write_satp = |_write_satp_T_14; // @[playground/src/pipeline/decode/Issue.scala 63:14]
  wire  _ret_T_2 = _csr_conflict_T & io_decodeInst_0_op == 7'ha; // @[playground/src/defines/Util.scala 14:31]
  wire  _ret_T_5 = _csr_conflict_T & io_decodeInst_0_op == 7'hb; // @[playground/src/defines/Util.scala 20:31]
  wire  _ret_T_6 = _ret_T_2 | _ret_T_5; // @[playground/src/defines/Util.scala 26:18]
  wire  _ret_T_9 = _csr_conflict_T_1 & io_decodeInst_1_op == 7'ha; // @[playground/src/defines/Util.scala 14:31]
  wire  _ret_T_12 = _csr_conflict_T_1 & io_decodeInst_1_op == 7'hb; // @[playground/src/defines/Util.scala 20:31]
  wire  _ret_T_13 = _ret_T_9 | _ret_T_12; // @[playground/src/defines/Util.scala 26:18]
  wire  ret = _ret_T_6 | _ret_T_13; // @[playground/src/pipeline/decode/Issue.scala 66:31]
  wire  is_some_csr_inst = write_satp | ret; // @[playground/src/pipeline/decode/Issue.scala 69:39]
  wire  single_issue = is_mou | is_bru | is_some_csr_inst; // @[playground/src/pipeline/decode/Issue.scala 72:41]
  wire  _io_inst1_allow_to_go_T = ~instFifo_invalid; // @[playground/src/pipeline/decode/Issue.scala 77:7]
  wire  _io_inst1_allow_to_go_T_1 = io_allow_to_go & _io_inst1_allow_to_go_T; // @[playground/src/pipeline/decode/Issue.scala 76:22]
  wire  _io_inst1_allow_to_go_T_2 = ~struct_conflict; // @[playground/src/pipeline/decode/Issue.scala 78:7]
  wire  _io_inst1_allow_to_go_T_3 = _io_inst1_allow_to_go_T_1 & _io_inst1_allow_to_go_T_2; // @[playground/src/pipeline/decode/Issue.scala 77:25]
  wire  _io_inst1_allow_to_go_T_4 = ~data_conflict; // @[playground/src/pipeline/decode/Issue.scala 79:7]
  wire  _io_inst1_allow_to_go_T_5 = _io_inst1_allow_to_go_T_3 & _io_inst1_allow_to_go_T_4; // @[playground/src/pipeline/decode/Issue.scala 78:24]
  wire  _io_inst1_allow_to_go_T_6 = ~single_issue; // @[playground/src/pipeline/decode/Issue.scala 80:7]
  assign io_inst1_allow_to_go = _io_inst1_allow_to_go_T_5 & _io_inst1_allow_to_go_T_6; // @[playground/src/pipeline/decode/Issue.scala 79:22]
endmodule
module DecodeUnit(
  output        io_instFifo_allow_to_go_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_instFifo_allow_to_go_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_instFifo_inst_0_inst, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [5:0]  io_instFifo_inst_0_pht_index, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_inst_0_addr_misaligned, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_inst_0_access_fault, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_inst_0_page_fault, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_instFifo_inst_0_pc, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_instFifo_inst_1_inst, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_inst_1_addr_misaligned, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_inst_1_access_fault, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_inst_1_page_fault, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_instFifo_inst_1_pc, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_info_empty, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_instFifo_info_almost_empty, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_regfile_0_src1_raddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_regfile_0_src1_rdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_regfile_0_src2_raddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_regfile_0_src2_rdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_regfile_1_src1_raddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_regfile_1_src1_rdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_regfile_1_src2_raddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_regfile_1_src2_rdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_forward_0_exe_wen, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [4:0]  io_forward_0_exe_waddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_forward_0_exe_wdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_forward_0_is_load, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_forward_0_mem_wen, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [4:0]  io_forward_0_mem_waddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_forward_0_mem_wdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_forward_1_exe_wen, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [4:0]  io_forward_1_exe_waddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_forward_1_exe_wdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_forward_1_is_load, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_forward_1_mem_wen, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [4:0]  io_forward_1_mem_waddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_forward_1_mem_wdata, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [1:0]  io_csr_mode, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [11:0] io_csr_interrupt, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_fetchUnit_branch, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_fetchUnit_target, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_bpu_pc, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_bpu_info_valid, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [2:0]  io_bpu_info_fusel, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [6:0]  io_bpu_info_op, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_bpu_info_imm, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [5:0]  io_bpu_pht_index, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_bpu_branch_inst, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_bpu_branch, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [63:0] io_bpu_target, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input  [5:0]  io_bpu_update_pht_index, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_pc, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_info_valid, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [2:0]  io_executeStage_inst_0_info_fusel, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [6:0]  io_executeStage_inst_0_info_op, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_info_reg_wen, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_executeStage_inst_0_info_reg_waddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_info_imm, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_info_inst, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_src_info_src1_data, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_src_info_src2_data, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_2, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_3, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_8, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_9, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_11, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_exception_12, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_2, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_3, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_4, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_5, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_6, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_7, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_8, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_9, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_10, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_0_ex_interrupt_11, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_ex_tval_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_ex_tval_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_ex_tval_2, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_0_ex_tval_12, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_pc, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_info_valid, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [2:0]  io_executeStage_inst_1_info_fusel, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [6:0]  io_executeStage_inst_1_info_op, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_info_reg_wen, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_executeStage_inst_1_info_reg_waddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_info_imm, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_info_inst, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_src_info_src1_data, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_src_info_src2_data, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_2, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_3, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_8, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_9, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_11, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_exception_12, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_2, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_3, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_4, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_5, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_6, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_7, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_8, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_9, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_10, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_inst_1_ex_interrupt_11, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_ex_tval_0, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_ex_tval_1, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_ex_tval_2, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_inst_1_ex_tval_12, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_jump_branch_info_jump_regiser, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_jump_branch_info_branch_inst, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_executeStage_jump_branch_info_pred_branch, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_jump_branch_info_branch_target, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [63:0] io_executeStage_jump_branch_info_update_pht_index, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_ctrl_inst0_src1_ren, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_ctrl_inst0_src1_raddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_ctrl_inst0_src2_ren, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output [4:0]  io_ctrl_inst0_src2_raddr, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  output        io_ctrl_branch, // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
  input         io_ctrl_allow_to_go // @[playground/src/pipeline/decode/DecodeUnit.scala 41:14]
);
  wire [63:0] decoder_0_io_in_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_0_io_out_info_inst_legal; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_0_io_out_info_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [4:0] decoder_0_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_0_io_out_info_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [4:0] decoder_0_io_out_info_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [2:0] decoder_0_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [6:0] decoder_0_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_0_io_out_info_reg_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [4:0] decoder_0_io_out_info_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [63:0] decoder_0_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [63:0] decoder_0_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [63:0] decoder_1_io_in_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_1_io_out_info_inst_legal; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_1_io_out_info_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [4:0] decoder_1_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_1_io_out_info_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [4:0] decoder_1_io_out_info_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [2:0] decoder_1_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [6:0] decoder_1_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  decoder_1_io_out_info_reg_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [4:0] decoder_1_io_out_info_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [63:0] decoder_1_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire [63:0] decoder_1_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
  wire  JumpCtrl_io_in_info_valid; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [4:0] JumpCtrl_io_in_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [2:0] JumpCtrl_io_in_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [6:0] JumpCtrl_io_in_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [63:0] JumpCtrl_io_in_src_info_src1_data; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [63:0] JumpCtrl_io_in_src_info_src2_data; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  JumpCtrl_io_in_forward_0_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [4:0] JumpCtrl_io_in_forward_0_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  JumpCtrl_io_in_forward_0_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [4:0] JumpCtrl_io_in_forward_0_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  JumpCtrl_io_in_forward_1_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [4:0] JumpCtrl_io_in_forward_1_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  JumpCtrl_io_in_forward_1_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [4:0] JumpCtrl_io_in_forward_1_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  JumpCtrl_io_out_jump_register; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  JumpCtrl_io_out_jump; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire [63:0] JumpCtrl_io_out_jump_target; // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
  wire  ForwardCtrl_io_in_forward_0_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_forward_0_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_forward_0_exe_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire  ForwardCtrl_io_in_forward_0_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire  ForwardCtrl_io_in_forward_0_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_forward_0_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_forward_0_mem_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire  ForwardCtrl_io_in_forward_1_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_forward_1_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_forward_1_exe_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire  ForwardCtrl_io_in_forward_1_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire  ForwardCtrl_io_in_forward_1_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_forward_1_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_forward_1_mem_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_regfile_0_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_regfile_0_src1_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_regfile_0_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_regfile_0_src2_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_regfile_1_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_regfile_1_src1_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [4:0] ForwardCtrl_io_in_regfile_1_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_in_regfile_1_src2_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_out_inst_0_src1_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_out_inst_0_src2_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_out_inst_1_src1_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire [63:0] ForwardCtrl_io_out_inst_1_src2_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
  wire  Issue_io_allow_to_go; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_instFifo_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_instFifo_almost_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [2:0] Issue_io_decodeInst_0_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [6:0] Issue_io_decodeInst_0_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_decodeInst_0_reg_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [4:0] Issue_io_decodeInst_0_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [63:0] Issue_io_decodeInst_0_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_decodeInst_1_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [4:0] Issue_io_decodeInst_1_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_decodeInst_1_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [4:0] Issue_io_decodeInst_1_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [2:0] Issue_io_decodeInst_1_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [6:0] Issue_io_decodeInst_1_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [63:0] Issue_io_decodeInst_1_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_execute_0_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [4:0] Issue_io_execute_0_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_execute_1_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire [4:0] Issue_io_execute_1_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  Issue_io_inst1_allow_to_go; // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
  wire  info_0_valid = ~io_instFifo_info_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 68:20]
  wire  inst0_branch = JumpCtrl_io_out_jump | io_bpu_branch; // @[playground/src/pipeline/decode/DecodeUnit.scala 90:40]
  wire [63:0] info_0_inst = decoder_0_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  _io_executeStage_inst_0_src_info_src1_data_T_2 = info_0_inst[6:0] == 7'h37; // @[playground/src/pipeline/decode/DecodeUnit.scala 119:29]
  wire [63:0] _io_executeStage_inst_0_src_info_src1_data_T_3 = _io_executeStage_inst_0_src_info_src1_data_T_2 ? 64'h0 :
    io_instFifo_inst_0_pc; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  info_0_src1_ren = decoder_0_io_out_info_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  info_0_src2_ren = decoder_0_io_out_info_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire [63:0] info_0_imm = decoder_0_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  info_0_inst_legal = decoder_0_io_out_info_inst_legal; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  _io_executeStage_inst_0_ex_exception_0_T_2 = |io_fetchUnit_target[1:0] & io_fetchUnit_branch; // @[playground/src/pipeline/decode/DecodeUnit.scala 133:60]
  wire [6:0] info_0_op = decoder_0_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire [2:0] info_0_fusel = decoder_0_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  _io_executeStage_inst_0_ex_exception_3_T_1 = info_0_fusel == 3'h3; // @[playground/src/pipeline/decode/DecodeUnit.scala 135:56]
  wire  _io_executeStage_inst_0_ex_exception_11_T = info_0_op == 7'h8; // @[playground/src/pipeline/decode/DecodeUnit.scala 137:18]
  wire [63:0] info_1_inst = decoder_1_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  _io_executeStage_inst_1_src_info_src1_data_T_2 = info_1_inst[6:0] == 7'h37; // @[playground/src/pipeline/decode/DecodeUnit.scala 119:29]
  wire [63:0] _io_executeStage_inst_1_src_info_src1_data_T_3 = _io_executeStage_inst_1_src_info_src1_data_T_2 ? 64'h0 :
    io_instFifo_inst_1_pc; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  info_1_src1_ren = decoder_1_io_out_info_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  info_1_src2_ren = decoder_1_io_out_info_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire [63:0] info_1_imm = decoder_1_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  info_1_inst_legal = decoder_1_io_out_info_inst_legal; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire [6:0] info_1_op = decoder_1_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire [2:0] info_1_fusel = decoder_1_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  wire  _io_executeStage_inst_1_ex_exception_3_T_1 = info_1_fusel == 3'h3; // @[playground/src/pipeline/decode/DecodeUnit.scala 135:56]
  wire  _io_executeStage_inst_1_ex_exception_11_T = info_1_op == 7'h8; // @[playground/src/pipeline/decode/DecodeUnit.scala 137:18]
  Decoder decoder_0 ( // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
    .io_in_inst(decoder_0_io_in_inst),
    .io_out_info_inst_legal(decoder_0_io_out_info_inst_legal),
    .io_out_info_src1_ren(decoder_0_io_out_info_src1_ren),
    .io_out_info_src1_raddr(decoder_0_io_out_info_src1_raddr),
    .io_out_info_src2_ren(decoder_0_io_out_info_src2_ren),
    .io_out_info_src2_raddr(decoder_0_io_out_info_src2_raddr),
    .io_out_info_fusel(decoder_0_io_out_info_fusel),
    .io_out_info_op(decoder_0_io_out_info_op),
    .io_out_info_reg_wen(decoder_0_io_out_info_reg_wen),
    .io_out_info_reg_waddr(decoder_0_io_out_info_reg_waddr),
    .io_out_info_imm(decoder_0_io_out_info_imm),
    .io_out_info_inst(decoder_0_io_out_info_inst)
  );
  Decoder decoder_1 ( // @[playground/src/pipeline/decode/DecodeUnit.scala 57:58]
    .io_in_inst(decoder_1_io_in_inst),
    .io_out_info_inst_legal(decoder_1_io_out_info_inst_legal),
    .io_out_info_src1_ren(decoder_1_io_out_info_src1_ren),
    .io_out_info_src1_raddr(decoder_1_io_out_info_src1_raddr),
    .io_out_info_src2_ren(decoder_1_io_out_info_src2_ren),
    .io_out_info_src2_raddr(decoder_1_io_out_info_src2_raddr),
    .io_out_info_fusel(decoder_1_io_out_info_fusel),
    .io_out_info_op(decoder_1_io_out_info_op),
    .io_out_info_reg_wen(decoder_1_io_out_info_reg_wen),
    .io_out_info_reg_waddr(decoder_1_io_out_info_reg_waddr),
    .io_out_info_imm(decoder_1_io_out_info_imm),
    .io_out_info_inst(decoder_1_io_out_info_inst)
  );
  JumpCtrl JumpCtrl ( // @[playground/src/pipeline/decode/DecodeUnit.scala 58:27]
    .io_in_info_valid(JumpCtrl_io_in_info_valid),
    .io_in_info_src1_raddr(JumpCtrl_io_in_info_src1_raddr),
    .io_in_info_fusel(JumpCtrl_io_in_info_fusel),
    .io_in_info_op(JumpCtrl_io_in_info_op),
    .io_in_src_info_src1_data(JumpCtrl_io_in_src_info_src1_data),
    .io_in_src_info_src2_data(JumpCtrl_io_in_src_info_src2_data),
    .io_in_forward_0_exe_wen(JumpCtrl_io_in_forward_0_exe_wen),
    .io_in_forward_0_exe_waddr(JumpCtrl_io_in_forward_0_exe_waddr),
    .io_in_forward_0_mem_wen(JumpCtrl_io_in_forward_0_mem_wen),
    .io_in_forward_0_mem_waddr(JumpCtrl_io_in_forward_0_mem_waddr),
    .io_in_forward_1_exe_wen(JumpCtrl_io_in_forward_1_exe_wen),
    .io_in_forward_1_exe_waddr(JumpCtrl_io_in_forward_1_exe_waddr),
    .io_in_forward_1_mem_wen(JumpCtrl_io_in_forward_1_mem_wen),
    .io_in_forward_1_mem_waddr(JumpCtrl_io_in_forward_1_mem_waddr),
    .io_out_jump_register(JumpCtrl_io_out_jump_register),
    .io_out_jump(JumpCtrl_io_out_jump),
    .io_out_jump_target(JumpCtrl_io_out_jump_target)
  );
  ForwardCtrl ForwardCtrl ( // @[playground/src/pipeline/decode/DecodeUnit.scala 59:27]
    .io_in_forward_0_exe_wen(ForwardCtrl_io_in_forward_0_exe_wen),
    .io_in_forward_0_exe_waddr(ForwardCtrl_io_in_forward_0_exe_waddr),
    .io_in_forward_0_exe_wdata(ForwardCtrl_io_in_forward_0_exe_wdata),
    .io_in_forward_0_is_load(ForwardCtrl_io_in_forward_0_is_load),
    .io_in_forward_0_mem_wen(ForwardCtrl_io_in_forward_0_mem_wen),
    .io_in_forward_0_mem_waddr(ForwardCtrl_io_in_forward_0_mem_waddr),
    .io_in_forward_0_mem_wdata(ForwardCtrl_io_in_forward_0_mem_wdata),
    .io_in_forward_1_exe_wen(ForwardCtrl_io_in_forward_1_exe_wen),
    .io_in_forward_1_exe_waddr(ForwardCtrl_io_in_forward_1_exe_waddr),
    .io_in_forward_1_exe_wdata(ForwardCtrl_io_in_forward_1_exe_wdata),
    .io_in_forward_1_is_load(ForwardCtrl_io_in_forward_1_is_load),
    .io_in_forward_1_mem_wen(ForwardCtrl_io_in_forward_1_mem_wen),
    .io_in_forward_1_mem_waddr(ForwardCtrl_io_in_forward_1_mem_waddr),
    .io_in_forward_1_mem_wdata(ForwardCtrl_io_in_forward_1_mem_wdata),
    .io_in_regfile_0_src1_raddr(ForwardCtrl_io_in_regfile_0_src1_raddr),
    .io_in_regfile_0_src1_rdata(ForwardCtrl_io_in_regfile_0_src1_rdata),
    .io_in_regfile_0_src2_raddr(ForwardCtrl_io_in_regfile_0_src2_raddr),
    .io_in_regfile_0_src2_rdata(ForwardCtrl_io_in_regfile_0_src2_rdata),
    .io_in_regfile_1_src1_raddr(ForwardCtrl_io_in_regfile_1_src1_raddr),
    .io_in_regfile_1_src1_rdata(ForwardCtrl_io_in_regfile_1_src1_rdata),
    .io_in_regfile_1_src2_raddr(ForwardCtrl_io_in_regfile_1_src2_raddr),
    .io_in_regfile_1_src2_rdata(ForwardCtrl_io_in_regfile_1_src2_rdata),
    .io_out_inst_0_src1_rdata(ForwardCtrl_io_out_inst_0_src1_rdata),
    .io_out_inst_0_src2_rdata(ForwardCtrl_io_out_inst_0_src2_rdata),
    .io_out_inst_1_src1_rdata(ForwardCtrl_io_out_inst_1_src1_rdata),
    .io_out_inst_1_src2_rdata(ForwardCtrl_io_out_inst_1_src2_rdata)
  );
  Issue Issue ( // @[playground/src/pipeline/decode/DecodeUnit.scala 60:27]
    .io_allow_to_go(Issue_io_allow_to_go),
    .io_instFifo_empty(Issue_io_instFifo_empty),
    .io_instFifo_almost_empty(Issue_io_instFifo_almost_empty),
    .io_decodeInst_0_fusel(Issue_io_decodeInst_0_fusel),
    .io_decodeInst_0_op(Issue_io_decodeInst_0_op),
    .io_decodeInst_0_reg_wen(Issue_io_decodeInst_0_reg_wen),
    .io_decodeInst_0_reg_waddr(Issue_io_decodeInst_0_reg_waddr),
    .io_decodeInst_0_inst(Issue_io_decodeInst_0_inst),
    .io_decodeInst_1_src1_ren(Issue_io_decodeInst_1_src1_ren),
    .io_decodeInst_1_src1_raddr(Issue_io_decodeInst_1_src1_raddr),
    .io_decodeInst_1_src2_ren(Issue_io_decodeInst_1_src2_ren),
    .io_decodeInst_1_src2_raddr(Issue_io_decodeInst_1_src2_raddr),
    .io_decodeInst_1_fusel(Issue_io_decodeInst_1_fusel),
    .io_decodeInst_1_op(Issue_io_decodeInst_1_op),
    .io_decodeInst_1_inst(Issue_io_decodeInst_1_inst),
    .io_execute_0_is_load(Issue_io_execute_0_is_load),
    .io_execute_0_reg_waddr(Issue_io_execute_0_reg_waddr),
    .io_execute_1_is_load(Issue_io_execute_1_is_load),
    .io_execute_1_reg_waddr(Issue_io_execute_1_reg_waddr),
    .io_inst1_allow_to_go(Issue_io_inst1_allow_to_go)
  );
  assign io_instFifo_allow_to_go_0 = io_ctrl_allow_to_go; // @[playground/src/pipeline/decode/DecodeUnit.scala 95:30]
  assign io_instFifo_allow_to_go_1 = Issue_io_inst1_allow_to_go; // @[playground/src/pipeline/decode/DecodeUnit.scala 73:30]
  assign io_regfile_0_src1_raddr = decoder_0_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_regfile_0_src2_raddr = decoder_0_io_out_info_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_regfile_1_src1_raddr = decoder_1_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_regfile_1_src2_raddr = decoder_1_io_out_info_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_fetchUnit_branch = inst0_branch & io_ctrl_allow_to_go; // @[playground/src/pipeline/decode/DecodeUnit.scala 92:39]
  assign io_fetchUnit_target = io_bpu_branch ? io_bpu_target : JumpCtrl_io_out_jump_target; // @[playground/src/pipeline/decode/DecodeUnit.scala 93:29]
  assign io_bpu_pc = io_instFifo_inst_0_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 96:30]
  assign io_bpu_info_valid = ~io_instFifo_info_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 68:20]
  assign io_bpu_info_fusel = decoder_0_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_bpu_info_op = decoder_0_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_bpu_info_imm = decoder_0_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_bpu_pht_index = io_instFifo_inst_0_pht_index; // @[playground/src/pipeline/decode/DecodeUnit.scala 98:30]
  assign io_executeStage_inst_0_pc = io_instFifo_inst_0_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 113:34]
  assign io_executeStage_inst_0_info_valid = ~io_instFifo_info_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 68:20]
  assign io_executeStage_inst_0_info_fusel = decoder_0_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_info_op = decoder_0_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_info_reg_wen = decoder_0_io_out_info_reg_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_info_reg_waddr = decoder_0_io_out_info_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_info_imm = decoder_0_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_info_inst = decoder_0_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_src_info_src1_data = info_0_src1_ren ? ForwardCtrl_io_out_inst_0_src1_rdata :
    _io_executeStage_inst_0_src_info_src1_data_T_3; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_executeStage_inst_0_src_info_src2_data = info_0_src2_ren ? ForwardCtrl_io_out_inst_0_src2_rdata : info_0_imm
    ; // @[playground/src/pipeline/decode/DecodeUnit.scala 122:54]
  assign io_executeStage_inst_0_ex_exception_0 = io_instFifo_inst_0_addr_misaligned |
    _io_executeStage_inst_0_ex_exception_0_T_2; // @[playground/src/pipeline/decode/DecodeUnit.scala 132:101]
  assign io_executeStage_inst_0_ex_exception_1 = io_instFifo_inst_0_access_fault; // @[playground/src/pipeline/decode/DecodeUnit.scala 130:59]
  assign io_executeStage_inst_0_ex_exception_2 = ~info_0_inst_legal; // @[playground/src/pipeline/decode/DecodeUnit.scala 129:62]
  assign io_executeStage_inst_0_ex_exception_3 = info_0_op == 7'h9 & info_0_fusel == 3'h3; // @[playground/src/pipeline/decode/DecodeUnit.scala 135:39]
  assign io_executeStage_inst_0_ex_exception_8 = _io_executeStage_inst_0_ex_exception_11_T & io_csr_mode == 2'h0 &
    _io_executeStage_inst_0_ex_exception_3_T_1; // @[playground/src/pipeline/decode/DecodeUnit.scala 141:56]
  assign io_executeStage_inst_0_ex_exception_9 = _io_executeStage_inst_0_ex_exception_11_T & io_csr_mode == 2'h1 &
    _io_executeStage_inst_0_ex_exception_3_T_1; // @[playground/src/pipeline/decode/DecodeUnit.scala 139:56]
  assign io_executeStage_inst_0_ex_exception_11 = info_0_op == 7'h8 & io_csr_mode == 2'h3 &
    _io_executeStage_inst_0_ex_exception_3_T_1; // @[playground/src/pipeline/decode/DecodeUnit.scala 137:56]
  assign io_executeStage_inst_0_ex_exception_12 = io_instFifo_inst_0_page_fault; // @[playground/src/pipeline/decode/DecodeUnit.scala 131:59]
  assign io_executeStage_inst_0_ex_interrupt_0 = io_csr_interrupt[0]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_1 = io_csr_interrupt[1]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_2 = io_csr_interrupt[2]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_3 = io_csr_interrupt[3]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_4 = io_csr_interrupt[4]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_5 = io_csr_interrupt[5]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_6 = io_csr_interrupt[6]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_7 = io_csr_interrupt[7]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_8 = io_csr_interrupt[8]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_9 = io_csr_interrupt[9]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_10 = io_csr_interrupt[10]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_interrupt_11 = io_csr_interrupt[11]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_0_ex_tval_0 = _io_executeStage_inst_0_ex_exception_0_T_2 ? io_fetchUnit_target :
    io_instFifo_inst_0_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 146:63]
  assign io_executeStage_inst_0_ex_tval_1 = io_instFifo_inst_0_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 144:54]
  assign io_executeStage_inst_0_ex_tval_2 = decoder_0_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_0_ex_tval_12 = io_instFifo_inst_0_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 143:54]
  assign io_executeStage_inst_1_pc = io_instFifo_inst_1_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 113:34]
  assign io_executeStage_inst_1_info_valid = ~io_instFifo_info_almost_empty & info_0_valid; // @[playground/src/pipeline/decode/DecodeUnit.scala 69:51]
  assign io_executeStage_inst_1_info_fusel = decoder_1_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_info_op = decoder_1_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_info_reg_wen = decoder_1_io_out_info_reg_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_info_reg_waddr = decoder_1_io_out_info_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_info_imm = decoder_1_io_out_info_imm; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_info_inst = decoder_1_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_src_info_src1_data = info_1_src1_ren ? ForwardCtrl_io_out_inst_1_src1_rdata :
    _io_executeStage_inst_1_src_info_src1_data_T_3; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_executeStage_inst_1_src_info_src2_data = info_1_src2_ren ? ForwardCtrl_io_out_inst_1_src2_rdata : info_1_imm
    ; // @[playground/src/pipeline/decode/DecodeUnit.scala 122:54]
  assign io_executeStage_inst_1_ex_exception_0 = io_instFifo_inst_1_addr_misaligned |
    _io_executeStage_inst_0_ex_exception_0_T_2; // @[playground/src/pipeline/decode/DecodeUnit.scala 132:101]
  assign io_executeStage_inst_1_ex_exception_1 = io_instFifo_inst_1_access_fault; // @[playground/src/pipeline/decode/DecodeUnit.scala 130:59]
  assign io_executeStage_inst_1_ex_exception_2 = ~info_1_inst_legal; // @[playground/src/pipeline/decode/DecodeUnit.scala 129:62]
  assign io_executeStage_inst_1_ex_exception_3 = info_1_op == 7'h9 & info_1_fusel == 3'h3; // @[playground/src/pipeline/decode/DecodeUnit.scala 135:39]
  assign io_executeStage_inst_1_ex_exception_8 = _io_executeStage_inst_1_ex_exception_11_T & io_csr_mode == 2'h0 &
    _io_executeStage_inst_1_ex_exception_3_T_1; // @[playground/src/pipeline/decode/DecodeUnit.scala 141:56]
  assign io_executeStage_inst_1_ex_exception_9 = _io_executeStage_inst_1_ex_exception_11_T & io_csr_mode == 2'h1 &
    _io_executeStage_inst_1_ex_exception_3_T_1; // @[playground/src/pipeline/decode/DecodeUnit.scala 139:56]
  assign io_executeStage_inst_1_ex_exception_11 = info_1_op == 7'h8 & io_csr_mode == 2'h3 &
    _io_executeStage_inst_1_ex_exception_3_T_1; // @[playground/src/pipeline/decode/DecodeUnit.scala 137:56]
  assign io_executeStage_inst_1_ex_exception_12 = io_instFifo_inst_1_page_fault; // @[playground/src/pipeline/decode/DecodeUnit.scala 131:59]
  assign io_executeStage_inst_1_ex_interrupt_0 = io_csr_interrupt[0]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_1 = io_csr_interrupt[1]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_2 = io_csr_interrupt[2]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_3 = io_csr_interrupt[3]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_4 = io_csr_interrupt[4]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_5 = io_csr_interrupt[5]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_6 = io_csr_interrupt[6]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_7 = io_csr_interrupt[7]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_8 = io_csr_interrupt[8]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_9 = io_csr_interrupt[9]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_10 = io_csr_interrupt[10]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_interrupt_11 = io_csr_interrupt[11]; // @[playground/src/pipeline/decode/DecodeUnit.scala 127:97]
  assign io_executeStage_inst_1_ex_tval_0 = _io_executeStage_inst_0_ex_exception_0_T_2 ? io_fetchUnit_target :
    io_instFifo_inst_1_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 146:63]
  assign io_executeStage_inst_1_ex_tval_1 = io_instFifo_inst_1_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 144:54]
  assign io_executeStage_inst_1_ex_tval_2 = decoder_1_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_executeStage_inst_1_ex_tval_12 = io_instFifo_inst_1_pc; // @[playground/src/pipeline/decode/DecodeUnit.scala 143:54]
  assign io_executeStage_jump_branch_info_jump_regiser = JumpCtrl_io_out_jump_register; // @[playground/src/pipeline/decode/DecodeUnit.scala 106:53]
  assign io_executeStage_jump_branch_info_branch_inst = io_bpu_branch_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 107:53]
  assign io_executeStage_jump_branch_info_pred_branch = io_bpu_branch; // @[playground/src/pipeline/decode/DecodeUnit.scala 108:53]
  assign io_executeStage_jump_branch_info_branch_target = io_bpu_target; // @[playground/src/pipeline/decode/DecodeUnit.scala 109:53]
  assign io_executeStage_jump_branch_info_update_pht_index = {{58'd0}, io_bpu_update_pht_index}; // @[playground/src/pipeline/decode/DecodeUnit.scala 110:53]
  assign io_ctrl_inst0_src1_ren = decoder_0_io_out_info_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_ctrl_inst0_src1_raddr = decoder_0_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_ctrl_inst0_src2_ren = decoder_0_io_out_info_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_ctrl_inst0_src2_raddr = decoder_0_io_out_info_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign io_ctrl_branch = io_fetchUnit_branch; // @[playground/src/pipeline/decode/DecodeUnit.scala 104:28]
  assign decoder_0_io_in_inst = io_instFifo_inst_0_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 75:32]
  assign decoder_1_io_in_inst = io_instFifo_inst_1_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 75:32]
  assign JumpCtrl_io_in_info_valid = ~io_instFifo_info_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 68:20]
  assign JumpCtrl_io_in_info_src1_raddr = decoder_0_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign JumpCtrl_io_in_info_fusel = decoder_0_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign JumpCtrl_io_in_info_op = decoder_0_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign JumpCtrl_io_in_src_info_src1_data = io_executeStage_inst_0_src_info_src1_data; // @[playground/src/pipeline/decode/DecodeUnit.scala 88:26]
  assign JumpCtrl_io_in_src_info_src2_data = io_executeStage_inst_0_src_info_src2_data; // @[playground/src/pipeline/decode/DecodeUnit.scala 88:26]
  assign JumpCtrl_io_in_forward_0_exe_wen = io_forward_0_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_0_exe_waddr = io_forward_0_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_0_mem_wen = io_forward_0_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_0_mem_waddr = io_forward_0_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_1_exe_wen = io_forward_1_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_1_exe_waddr = io_forward_1_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_1_mem_wen = io_forward_1_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign JumpCtrl_io_in_forward_1_mem_waddr = io_forward_1_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 86:26]
  assign ForwardCtrl_io_in_forward_0_exe_wen = io_forward_0_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_0_exe_waddr = io_forward_0_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_0_exe_wdata = io_forward_0_exe_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_0_is_load = io_forward_0_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_0_mem_wen = io_forward_0_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_0_mem_waddr = io_forward_0_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_0_mem_wdata = io_forward_0_mem_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_exe_wen = io_forward_1_exe_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_exe_waddr = io_forward_1_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_exe_wdata = io_forward_1_exe_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_is_load = io_forward_1_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_mem_wen = io_forward_1_mem_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_mem_waddr = io_forward_1_mem_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_forward_1_mem_wdata = io_forward_1_mem_wdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 83:26]
  assign ForwardCtrl_io_in_regfile_0_src1_raddr = io_regfile_0_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_0_src1_rdata = io_regfile_0_src1_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_0_src2_raddr = io_regfile_0_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_0_src2_rdata = io_regfile_0_src2_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_1_src1_raddr = io_regfile_1_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_1_src1_rdata = io_regfile_1_src1_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_1_src2_raddr = io_regfile_1_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign ForwardCtrl_io_in_regfile_1_src2_rdata = io_regfile_1_src2_rdata; // @[playground/src/pipeline/decode/DecodeUnit.scala 84:26]
  assign Issue_io_allow_to_go = io_ctrl_allow_to_go; // @[playground/src/pipeline/decode/DecodeUnit.scala 71:30]
  assign Issue_io_instFifo_empty = io_instFifo_info_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 72:30]
  assign Issue_io_instFifo_almost_empty = io_instFifo_info_almost_empty; // @[playground/src/pipeline/decode/DecodeUnit.scala 72:30]
  assign Issue_io_decodeInst_0_fusel = decoder_0_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_0_op = decoder_0_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_0_reg_wen = decoder_0_io_out_info_reg_wen; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_0_reg_waddr = decoder_0_io_out_info_reg_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_0_inst = decoder_0_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_src1_ren = decoder_1_io_out_info_src1_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_src1_raddr = decoder_1_io_out_info_src1_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_src2_ren = decoder_1_io_out_info_src2_ren; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_src2_raddr = decoder_1_io_out_info_src2_raddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_fusel = decoder_1_io_out_info_fusel; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_op = decoder_1_io_out_info_op; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_decodeInst_1_inst = decoder_1_io_out_info_inst; // @[playground/src/pipeline/decode/DecodeUnit.scala 64:18 67:17]
  assign Issue_io_execute_0_is_load = io_forward_0_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 77:32]
  assign Issue_io_execute_0_reg_waddr = io_forward_0_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 78:32]
  assign Issue_io_execute_1_is_load = io_forward_1_is_load; // @[playground/src/pipeline/decode/DecodeUnit.scala 77:32]
  assign Issue_io_execute_1_reg_waddr = io_forward_1_exe_waddr; // @[playground/src/pipeline/decode/DecodeUnit.scala 78:32]
endmodule
module ARegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_read_0_src1_raddr, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  output [63:0] io_read_0_src1_rdata, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [4:0]  io_read_0_src2_raddr, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  output [63:0] io_read_0_src2_rdata, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [4:0]  io_read_1_src1_raddr, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  output [63:0] io_read_1_src1_rdata, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [4:0]  io_read_1_src2_raddr, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  output [63:0] io_read_1_src2_rdata, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input         io_write_0_wen, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [4:0]  io_write_0_waddr, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [63:0] io_write_0_wdata, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input         io_write_1_wen, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [4:0]  io_write_1_waddr, // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
  input  [63:0] io_write_1_wdata // @[playground/src/pipeline/decode/ARegfile.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_1; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_2; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_3; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_4; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_5; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_6; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_7; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_8; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_9; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_10; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_11; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_12; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_13; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_14; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_15; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_16; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_17; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_18; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_19; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_20; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_21; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_22; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_23; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_24; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_25; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_26; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_27; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_28; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_29; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_30; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  reg [63:0] regs_31; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
  wire [63:0] _GEN_0 = 5'h0 == io_write_0_waddr ? io_write_0_wdata : regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_1 = 5'h1 == io_write_0_waddr ? io_write_0_wdata : regs_1; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_2 = 5'h2 == io_write_0_waddr ? io_write_0_wdata : regs_2; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_3 = 5'h3 == io_write_0_waddr ? io_write_0_wdata : regs_3; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_4 = 5'h4 == io_write_0_waddr ? io_write_0_wdata : regs_4; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_5 = 5'h5 == io_write_0_waddr ? io_write_0_wdata : regs_5; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_6 = 5'h6 == io_write_0_waddr ? io_write_0_wdata : regs_6; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_7 = 5'h7 == io_write_0_waddr ? io_write_0_wdata : regs_7; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_8 = 5'h8 == io_write_0_waddr ? io_write_0_wdata : regs_8; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_9 = 5'h9 == io_write_0_waddr ? io_write_0_wdata : regs_9; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_10 = 5'ha == io_write_0_waddr ? io_write_0_wdata : regs_10; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_11 = 5'hb == io_write_0_waddr ? io_write_0_wdata : regs_11; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_12 = 5'hc == io_write_0_waddr ? io_write_0_wdata : regs_12; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_13 = 5'hd == io_write_0_waddr ? io_write_0_wdata : regs_13; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_14 = 5'he == io_write_0_waddr ? io_write_0_wdata : regs_14; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_15 = 5'hf == io_write_0_waddr ? io_write_0_wdata : regs_15; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_16 = 5'h10 == io_write_0_waddr ? io_write_0_wdata : regs_16; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_17 = 5'h11 == io_write_0_waddr ? io_write_0_wdata : regs_17; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_18 = 5'h12 == io_write_0_waddr ? io_write_0_wdata : regs_18; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_19 = 5'h13 == io_write_0_waddr ? io_write_0_wdata : regs_19; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_20 = 5'h14 == io_write_0_waddr ? io_write_0_wdata : regs_20; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_21 = 5'h15 == io_write_0_waddr ? io_write_0_wdata : regs_21; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_22 = 5'h16 == io_write_0_waddr ? io_write_0_wdata : regs_22; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_23 = 5'h17 == io_write_0_waddr ? io_write_0_wdata : regs_23; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_24 = 5'h18 == io_write_0_waddr ? io_write_0_wdata : regs_24; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_25 = 5'h19 == io_write_0_waddr ? io_write_0_wdata : regs_25; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_26 = 5'h1a == io_write_0_waddr ? io_write_0_wdata : regs_26; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_27 = 5'h1b == io_write_0_waddr ? io_write_0_wdata : regs_27; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_28 = 5'h1c == io_write_0_waddr ? io_write_0_wdata : regs_28; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_29 = 5'h1d == io_write_0_waddr ? io_write_0_wdata : regs_29; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_30 = 5'h1e == io_write_0_waddr ? io_write_0_wdata : regs_30; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_31 = 5'h1f == io_write_0_waddr ? io_write_0_wdata : regs_31; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 37:{31,31}]
  wire [63:0] _GEN_32 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_0 : regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_33 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_1 : regs_1; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_34 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_2 : regs_2; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_35 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_3 : regs_3; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_36 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_4 : regs_4; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_37 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_5 : regs_5; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_38 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_6 : regs_6; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_39 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_7 : regs_7; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_40 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_8 : regs_8; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_41 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_9 : regs_9; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_42 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_10 : regs_10; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_43 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_11 : regs_11; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_44 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_12 : regs_12; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_45 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_13 : regs_13; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_46 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_14 : regs_14; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_47 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_15 : regs_15; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_48 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_16 : regs_16; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_49 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_17 : regs_17; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_50 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_18 : regs_18; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_51 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_19 : regs_19; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_52 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_20 : regs_20; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_53 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_21 : regs_21; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_54 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_22 : regs_22; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_55 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_23 : regs_23; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_56 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_24 : regs_24; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_57 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_25 : regs_25; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_58 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_26 : regs_26; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_59 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_27 : regs_27; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_60 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_28 : regs_28; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_61 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_29 : regs_29; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_62 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_30 : regs_30; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_63 = io_write_0_wen & io_write_0_waddr != 5'h0 ? _GEN_31 : regs_31; // @[playground/src/pipeline/decode/ARegfile.scala 32:21 36:56]
  wire [63:0] _GEN_129 = 5'h1 == io_read_0_src1_raddr ? regs_1 : regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_130 = 5'h2 == io_read_0_src1_raddr ? regs_2 : _GEN_129; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_131 = 5'h3 == io_read_0_src1_raddr ? regs_3 : _GEN_130; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_132 = 5'h4 == io_read_0_src1_raddr ? regs_4 : _GEN_131; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_133 = 5'h5 == io_read_0_src1_raddr ? regs_5 : _GEN_132; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_134 = 5'h6 == io_read_0_src1_raddr ? regs_6 : _GEN_133; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_135 = 5'h7 == io_read_0_src1_raddr ? regs_7 : _GEN_134; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_136 = 5'h8 == io_read_0_src1_raddr ? regs_8 : _GEN_135; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_137 = 5'h9 == io_read_0_src1_raddr ? regs_9 : _GEN_136; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_138 = 5'ha == io_read_0_src1_raddr ? regs_10 : _GEN_137; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_139 = 5'hb == io_read_0_src1_raddr ? regs_11 : _GEN_138; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_140 = 5'hc == io_read_0_src1_raddr ? regs_12 : _GEN_139; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_141 = 5'hd == io_read_0_src1_raddr ? regs_13 : _GEN_140; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_142 = 5'he == io_read_0_src1_raddr ? regs_14 : _GEN_141; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_143 = 5'hf == io_read_0_src1_raddr ? regs_15 : _GEN_142; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_144 = 5'h10 == io_read_0_src1_raddr ? regs_16 : _GEN_143; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_145 = 5'h11 == io_read_0_src1_raddr ? regs_17 : _GEN_144; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_146 = 5'h12 == io_read_0_src1_raddr ? regs_18 : _GEN_145; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_147 = 5'h13 == io_read_0_src1_raddr ? regs_19 : _GEN_146; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_148 = 5'h14 == io_read_0_src1_raddr ? regs_20 : _GEN_147; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_149 = 5'h15 == io_read_0_src1_raddr ? regs_21 : _GEN_148; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_150 = 5'h16 == io_read_0_src1_raddr ? regs_22 : _GEN_149; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_151 = 5'h17 == io_read_0_src1_raddr ? regs_23 : _GEN_150; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_152 = 5'h18 == io_read_0_src1_raddr ? regs_24 : _GEN_151; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_153 = 5'h19 == io_read_0_src1_raddr ? regs_25 : _GEN_152; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_154 = 5'h1a == io_read_0_src1_raddr ? regs_26 : _GEN_153; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_155 = 5'h1b == io_read_0_src1_raddr ? regs_27 : _GEN_154; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_156 = 5'h1c == io_read_0_src1_raddr ? regs_28 : _GEN_155; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_157 = 5'h1d == io_read_0_src1_raddr ? regs_29 : _GEN_156; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_158 = 5'h1e == io_read_0_src1_raddr ? regs_30 : _GEN_157; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_159 = 5'h1f == io_read_0_src1_raddr ? regs_31 : _GEN_158; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_160 = io_write_0_wen & io_read_0_src1_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_159; // @[playground/src/pipeline/decode/ARegfile.scala 47:29 49:78 50:33]
  wire [63:0] _GEN_161 = io_write_1_wen & io_read_0_src1_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_160; // @[playground/src/pipeline/decode/ARegfile.scala 49:78 50:33]
  wire [63:0] _GEN_164 = 5'h1 == io_read_0_src2_raddr ? regs_1 : regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_165 = 5'h2 == io_read_0_src2_raddr ? regs_2 : _GEN_164; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_166 = 5'h3 == io_read_0_src2_raddr ? regs_3 : _GEN_165; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_167 = 5'h4 == io_read_0_src2_raddr ? regs_4 : _GEN_166; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_168 = 5'h5 == io_read_0_src2_raddr ? regs_5 : _GEN_167; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_169 = 5'h6 == io_read_0_src2_raddr ? regs_6 : _GEN_168; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_170 = 5'h7 == io_read_0_src2_raddr ? regs_7 : _GEN_169; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_171 = 5'h8 == io_read_0_src2_raddr ? regs_8 : _GEN_170; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_172 = 5'h9 == io_read_0_src2_raddr ? regs_9 : _GEN_171; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_173 = 5'ha == io_read_0_src2_raddr ? regs_10 : _GEN_172; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_174 = 5'hb == io_read_0_src2_raddr ? regs_11 : _GEN_173; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_175 = 5'hc == io_read_0_src2_raddr ? regs_12 : _GEN_174; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_176 = 5'hd == io_read_0_src2_raddr ? regs_13 : _GEN_175; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_177 = 5'he == io_read_0_src2_raddr ? regs_14 : _GEN_176; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_178 = 5'hf == io_read_0_src2_raddr ? regs_15 : _GEN_177; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_179 = 5'h10 == io_read_0_src2_raddr ? regs_16 : _GEN_178; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_180 = 5'h11 == io_read_0_src2_raddr ? regs_17 : _GEN_179; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_181 = 5'h12 == io_read_0_src2_raddr ? regs_18 : _GEN_180; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_182 = 5'h13 == io_read_0_src2_raddr ? regs_19 : _GEN_181; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_183 = 5'h14 == io_read_0_src2_raddr ? regs_20 : _GEN_182; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_184 = 5'h15 == io_read_0_src2_raddr ? regs_21 : _GEN_183; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_185 = 5'h16 == io_read_0_src2_raddr ? regs_22 : _GEN_184; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_186 = 5'h17 == io_read_0_src2_raddr ? regs_23 : _GEN_185; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_187 = 5'h18 == io_read_0_src2_raddr ? regs_24 : _GEN_186; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_188 = 5'h19 == io_read_0_src2_raddr ? regs_25 : _GEN_187; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_189 = 5'h1a == io_read_0_src2_raddr ? regs_26 : _GEN_188; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_190 = 5'h1b == io_read_0_src2_raddr ? regs_27 : _GEN_189; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_191 = 5'h1c == io_read_0_src2_raddr ? regs_28 : _GEN_190; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_192 = 5'h1d == io_read_0_src2_raddr ? regs_29 : _GEN_191; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_193 = 5'h1e == io_read_0_src2_raddr ? regs_30 : _GEN_192; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_194 = 5'h1f == io_read_0_src2_raddr ? regs_31 : _GEN_193; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_195 = io_write_0_wen & io_read_0_src2_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_194; // @[playground/src/pipeline/decode/ARegfile.scala 58:29 60:78 61:33]
  wire [63:0] _GEN_196 = io_write_1_wen & io_read_0_src2_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_195; // @[playground/src/pipeline/decode/ARegfile.scala 60:78 61:33]
  wire [63:0] _GEN_199 = 5'h1 == io_read_1_src1_raddr ? regs_1 : regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_200 = 5'h2 == io_read_1_src1_raddr ? regs_2 : _GEN_199; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_201 = 5'h3 == io_read_1_src1_raddr ? regs_3 : _GEN_200; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_202 = 5'h4 == io_read_1_src1_raddr ? regs_4 : _GEN_201; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_203 = 5'h5 == io_read_1_src1_raddr ? regs_5 : _GEN_202; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_204 = 5'h6 == io_read_1_src1_raddr ? regs_6 : _GEN_203; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_205 = 5'h7 == io_read_1_src1_raddr ? regs_7 : _GEN_204; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_206 = 5'h8 == io_read_1_src1_raddr ? regs_8 : _GEN_205; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_207 = 5'h9 == io_read_1_src1_raddr ? regs_9 : _GEN_206; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_208 = 5'ha == io_read_1_src1_raddr ? regs_10 : _GEN_207; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_209 = 5'hb == io_read_1_src1_raddr ? regs_11 : _GEN_208; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_210 = 5'hc == io_read_1_src1_raddr ? regs_12 : _GEN_209; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_211 = 5'hd == io_read_1_src1_raddr ? regs_13 : _GEN_210; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_212 = 5'he == io_read_1_src1_raddr ? regs_14 : _GEN_211; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_213 = 5'hf == io_read_1_src1_raddr ? regs_15 : _GEN_212; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_214 = 5'h10 == io_read_1_src1_raddr ? regs_16 : _GEN_213; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_215 = 5'h11 == io_read_1_src1_raddr ? regs_17 : _GEN_214; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_216 = 5'h12 == io_read_1_src1_raddr ? regs_18 : _GEN_215; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_217 = 5'h13 == io_read_1_src1_raddr ? regs_19 : _GEN_216; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_218 = 5'h14 == io_read_1_src1_raddr ? regs_20 : _GEN_217; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_219 = 5'h15 == io_read_1_src1_raddr ? regs_21 : _GEN_218; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_220 = 5'h16 == io_read_1_src1_raddr ? regs_22 : _GEN_219; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_221 = 5'h17 == io_read_1_src1_raddr ? regs_23 : _GEN_220; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_222 = 5'h18 == io_read_1_src1_raddr ? regs_24 : _GEN_221; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_223 = 5'h19 == io_read_1_src1_raddr ? regs_25 : _GEN_222; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_224 = 5'h1a == io_read_1_src1_raddr ? regs_26 : _GEN_223; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_225 = 5'h1b == io_read_1_src1_raddr ? regs_27 : _GEN_224; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_226 = 5'h1c == io_read_1_src1_raddr ? regs_28 : _GEN_225; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_227 = 5'h1d == io_read_1_src1_raddr ? regs_29 : _GEN_226; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_228 = 5'h1e == io_read_1_src1_raddr ? regs_30 : _GEN_227; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_229 = 5'h1f == io_read_1_src1_raddr ? regs_31 : _GEN_228; // @[playground/src/pipeline/decode/ARegfile.scala 47:{29,29}]
  wire [63:0] _GEN_230 = io_write_0_wen & io_read_1_src1_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_229; // @[playground/src/pipeline/decode/ARegfile.scala 47:29 49:78 50:33]
  wire [63:0] _GEN_231 = io_write_1_wen & io_read_1_src1_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_230; // @[playground/src/pipeline/decode/ARegfile.scala 49:78 50:33]
  wire [63:0] _GEN_234 = 5'h1 == io_read_1_src2_raddr ? regs_1 : regs_0; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_235 = 5'h2 == io_read_1_src2_raddr ? regs_2 : _GEN_234; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_236 = 5'h3 == io_read_1_src2_raddr ? regs_3 : _GEN_235; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_237 = 5'h4 == io_read_1_src2_raddr ? regs_4 : _GEN_236; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_238 = 5'h5 == io_read_1_src2_raddr ? regs_5 : _GEN_237; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_239 = 5'h6 == io_read_1_src2_raddr ? regs_6 : _GEN_238; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_240 = 5'h7 == io_read_1_src2_raddr ? regs_7 : _GEN_239; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_241 = 5'h8 == io_read_1_src2_raddr ? regs_8 : _GEN_240; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_242 = 5'h9 == io_read_1_src2_raddr ? regs_9 : _GEN_241; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_243 = 5'ha == io_read_1_src2_raddr ? regs_10 : _GEN_242; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_244 = 5'hb == io_read_1_src2_raddr ? regs_11 : _GEN_243; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_245 = 5'hc == io_read_1_src2_raddr ? regs_12 : _GEN_244; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_246 = 5'hd == io_read_1_src2_raddr ? regs_13 : _GEN_245; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_247 = 5'he == io_read_1_src2_raddr ? regs_14 : _GEN_246; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_248 = 5'hf == io_read_1_src2_raddr ? regs_15 : _GEN_247; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_249 = 5'h10 == io_read_1_src2_raddr ? regs_16 : _GEN_248; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_250 = 5'h11 == io_read_1_src2_raddr ? regs_17 : _GEN_249; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_251 = 5'h12 == io_read_1_src2_raddr ? regs_18 : _GEN_250; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_252 = 5'h13 == io_read_1_src2_raddr ? regs_19 : _GEN_251; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_253 = 5'h14 == io_read_1_src2_raddr ? regs_20 : _GEN_252; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_254 = 5'h15 == io_read_1_src2_raddr ? regs_21 : _GEN_253; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_255 = 5'h16 == io_read_1_src2_raddr ? regs_22 : _GEN_254; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_256 = 5'h17 == io_read_1_src2_raddr ? regs_23 : _GEN_255; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_257 = 5'h18 == io_read_1_src2_raddr ? regs_24 : _GEN_256; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_258 = 5'h19 == io_read_1_src2_raddr ? regs_25 : _GEN_257; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_259 = 5'h1a == io_read_1_src2_raddr ? regs_26 : _GEN_258; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_260 = 5'h1b == io_read_1_src2_raddr ? regs_27 : _GEN_259; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_261 = 5'h1c == io_read_1_src2_raddr ? regs_28 : _GEN_260; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_262 = 5'h1d == io_read_1_src2_raddr ? regs_29 : _GEN_261; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_263 = 5'h1e == io_read_1_src2_raddr ? regs_30 : _GEN_262; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_264 = 5'h1f == io_read_1_src2_raddr ? regs_31 : _GEN_263; // @[playground/src/pipeline/decode/ARegfile.scala 58:{29,29}]
  wire [63:0] _GEN_265 = io_write_0_wen & io_read_1_src2_raddr == io_write_0_waddr ? io_write_0_wdata : _GEN_264; // @[playground/src/pipeline/decode/ARegfile.scala 58:29 60:78 61:33]
  wire [63:0] _GEN_266 = io_write_1_wen & io_read_1_src2_raddr == io_write_1_waddr ? io_write_1_wdata : _GEN_265; // @[playground/src/pipeline/decode/ARegfile.scala 60:78 61:33]
  assign io_read_0_src1_rdata = io_read_0_src1_raddr == 5'h0 ? 64'h0 : _GEN_161; // @[playground/src/pipeline/decode/ARegfile.scala 44:41 45:29]
  assign io_read_0_src2_rdata = io_read_0_src2_raddr == 5'h0 ? 64'h0 : _GEN_196; // @[playground/src/pipeline/decode/ARegfile.scala 55:41 56:29]
  assign io_read_1_src1_rdata = io_read_1_src1_raddr == 5'h0 ? 64'h0 : _GEN_231; // @[playground/src/pipeline/decode/ARegfile.scala 44:41 45:29]
  assign io_read_1_src2_rdata = io_read_1_src2_raddr == 5'h0 ? 64'h0 : _GEN_266; // @[playground/src/pipeline/decode/ARegfile.scala 55:41 56:29]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_0 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h0 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_0 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_0 <= _GEN_32;
      end
    end else begin
      regs_0 <= _GEN_32;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_1 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_1 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_1 <= _GEN_33;
      end
    end else begin
      regs_1 <= _GEN_33;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_2 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h2 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_2 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_2 <= _GEN_34;
      end
    end else begin
      regs_2 <= _GEN_34;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_3 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h3 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_3 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_3 <= _GEN_35;
      end
    end else begin
      regs_3 <= _GEN_35;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_4 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h4 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_4 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_4 <= _GEN_36;
      end
    end else begin
      regs_4 <= _GEN_36;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_5 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h5 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_5 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_5 <= _GEN_37;
      end
    end else begin
      regs_5 <= _GEN_37;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_6 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h6 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_6 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_6 <= _GEN_38;
      end
    end else begin
      regs_6 <= _GEN_38;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_7 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h7 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_7 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_7 <= _GEN_39;
      end
    end else begin
      regs_7 <= _GEN_39;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_8 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h8 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_8 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_8 <= _GEN_40;
      end
    end else begin
      regs_8 <= _GEN_40;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_9 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h9 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_9 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_9 <= _GEN_41;
      end
    end else begin
      regs_9 <= _GEN_41;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_10 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'ha == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_10 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_10 <= _GEN_42;
      end
    end else begin
      regs_10 <= _GEN_42;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_11 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'hb == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_11 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_11 <= _GEN_43;
      end
    end else begin
      regs_11 <= _GEN_43;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_12 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'hc == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_12 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_12 <= _GEN_44;
      end
    end else begin
      regs_12 <= _GEN_44;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_13 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'hd == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_13 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_13 <= _GEN_45;
      end
    end else begin
      regs_13 <= _GEN_45;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_14 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'he == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_14 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_14 <= _GEN_46;
      end
    end else begin
      regs_14 <= _GEN_46;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_15 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'hf == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_15 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_15 <= _GEN_47;
      end
    end else begin
      regs_15 <= _GEN_47;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_16 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h10 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_16 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_16 <= _GEN_48;
      end
    end else begin
      regs_16 <= _GEN_48;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_17 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h11 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_17 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_17 <= _GEN_49;
      end
    end else begin
      regs_17 <= _GEN_49;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_18 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h12 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_18 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_18 <= _GEN_50;
      end
    end else begin
      regs_18 <= _GEN_50;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_19 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h13 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_19 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_19 <= _GEN_51;
      end
    end else begin
      regs_19 <= _GEN_51;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_20 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h14 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_20 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_20 <= _GEN_52;
      end
    end else begin
      regs_20 <= _GEN_52;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_21 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h15 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_21 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_21 <= _GEN_53;
      end
    end else begin
      regs_21 <= _GEN_53;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_22 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h16 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_22 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_22 <= _GEN_54;
      end
    end else begin
      regs_22 <= _GEN_54;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_23 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h17 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_23 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_23 <= _GEN_55;
      end
    end else begin
      regs_23 <= _GEN_55;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_24 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h18 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_24 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_24 <= _GEN_56;
      end
    end else begin
      regs_24 <= _GEN_56;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_25 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h19 == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_25 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_25 <= _GEN_57;
      end
    end else begin
      regs_25 <= _GEN_57;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_26 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1a == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_26 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_26 <= _GEN_58;
      end
    end else begin
      regs_26 <= _GEN_58;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_27 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1b == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_27 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_27 <= _GEN_59;
      end
    end else begin
      regs_27 <= _GEN_59;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_28 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1c == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_28 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_28 <= _GEN_60;
      end
    end else begin
      regs_28 <= _GEN_60;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_29 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1d == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_29 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_29 <= _GEN_61;
      end
    end else begin
      regs_29 <= _GEN_61;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_30 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1e == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_30 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_30 <= _GEN_62;
      end
    end else begin
      regs_30 <= _GEN_62;
    end
    if (reset) begin // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
      regs_31 <= 64'h0; // @[playground/src/pipeline/decode/ARegfile.scala 32:21]
    end else if (io_write_1_wen & io_write_1_waddr != 5'h0) begin // @[playground/src/pipeline/decode/ARegfile.scala 36:56]
      if (5'h1f == io_write_1_waddr) begin // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
        regs_31 <= io_write_1_wdata; // @[playground/src/pipeline/decode/ARegfile.scala 37:31]
      end else begin
        regs_31 <= _GEN_63;
      end
    end else begin
      regs_31 <= _GEN_63;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ExecuteStage(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_ctrl_allow_to_go_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_ctrl_clear_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_ctrl_clear_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_pc, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_info_valid, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [2:0]  io_decodeUnit_inst_0_info_fusel, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [6:0]  io_decodeUnit_inst_0_info_op, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [4:0]  io_decodeUnit_inst_0_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_info_imm, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_info_inst, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_0_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_0_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_pc, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_info_valid, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [2:0]  io_decodeUnit_inst_1_info_fusel, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [6:0]  io_decodeUnit_inst_1_info_op, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [4:0]  io_decodeUnit_inst_1_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_info_imm, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_info_inst, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_inst_1_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_inst_1_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_jump_branch_info_jump_regiser, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_jump_branch_info_branch_inst, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input         io_decodeUnit_jump_branch_info_pred_branch, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_jump_branch_info_branch_target, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  input  [63:0] io_decodeUnit_jump_branch_info_update_pht_index, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_pc, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_info_valid, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [2:0]  io_executeUnit_inst_0_info_fusel, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [6:0]  io_executeUnit_inst_0_info_op, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [4:0]  io_executeUnit_inst_0_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_info_imm, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_info_inst, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_0_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_0_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_pc, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_info_valid, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [2:0]  io_executeUnit_inst_1_info_fusel, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [6:0]  io_executeUnit_inst_1_info_op, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [4:0]  io_executeUnit_inst_1_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_info_imm, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_info_inst, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_inst_1_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_inst_1_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_jump_branch_info_jump_regiser, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_jump_branch_info_branch_inst, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output        io_executeUnit_jump_branch_info_pred_branch, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_jump_branch_info_branch_target, // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
  output [63:0] io_executeUnit_jump_branch_info_update_pht_index // @[playground/src/pipeline/execute/ExecuteStage.scala 31:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] inst_0_pc; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [2:0] inst_0_info_fusel; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [6:0] inst_0_info_op; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [4:0] inst_0_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_info_imm; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_info_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_0_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_ex_tval_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_0_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_pc; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [2:0] inst_1_info_fusel; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [6:0] inst_1_info_op; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [4:0] inst_1_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_info_imm; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_info_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  inst_1_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_ex_tval_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg [63:0] inst_1_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
  reg  jump_branch_info_jump_regiser; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
  reg  jump_branch_info_branch_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
  reg  jump_branch_info_pred_branch; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
  reg [63:0] jump_branch_info_branch_target; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
  reg [63:0] jump_branch_info_update_pht_index; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
  assign io_executeUnit_inst_0_pc = inst_0_pc; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_valid = inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_fusel = inst_0_info_fusel; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_op = inst_0_info_op; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_reg_wen = inst_0_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_reg_waddr = inst_0_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_imm = inst_0_info_imm; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_info_inst = inst_0_info_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_src_info_src1_data = inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_src_info_src2_data = inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_0 = inst_0_ex_exception_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_1 = inst_0_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_2 = inst_0_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_3 = inst_0_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_8 = inst_0_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_9 = inst_0_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_11 = inst_0_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_exception_12 = inst_0_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_0 = inst_0_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_1 = inst_0_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_2 = inst_0_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_3 = inst_0_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_4 = inst_0_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_5 = inst_0_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_6 = inst_0_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_7 = inst_0_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_8 = inst_0_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_9 = inst_0_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_10 = inst_0_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_interrupt_11 = inst_0_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_tval_0 = inst_0_ex_tval_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_tval_1 = inst_0_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_tval_2 = inst_0_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_0_ex_tval_12 = inst_0_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_pc = inst_1_pc; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_valid = inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_fusel = inst_1_info_fusel; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_op = inst_1_info_op; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_reg_wen = inst_1_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_reg_waddr = inst_1_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_imm = inst_1_info_imm; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_info_inst = inst_1_info_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_src_info_src1_data = inst_1_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_src_info_src2_data = inst_1_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_0 = inst_1_ex_exception_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_1 = inst_1_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_2 = inst_1_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_3 = inst_1_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_8 = inst_1_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_9 = inst_1_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_11 = inst_1_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_exception_12 = inst_1_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_0 = inst_1_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_1 = inst_1_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_2 = inst_1_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_3 = inst_1_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_4 = inst_1_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_5 = inst_1_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_6 = inst_1_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_7 = inst_1_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_8 = inst_1_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_9 = inst_1_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_10 = inst_1_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_interrupt_11 = inst_1_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_tval_0 = inst_1_ex_tval_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_tval_1 = inst_1_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_tval_2 = inst_1_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_inst_1_ex_tval_12 = inst_1_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 58:35]
  assign io_executeUnit_jump_branch_info_jump_regiser = jump_branch_info_jump_regiser; // @[playground/src/pipeline/execute/ExecuteStage.scala 59:35]
  assign io_executeUnit_jump_branch_info_branch_inst = jump_branch_info_branch_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 59:35]
  assign io_executeUnit_jump_branch_info_pred_branch = jump_branch_info_pred_branch; // @[playground/src/pipeline/execute/ExecuteStage.scala 59:35]
  assign io_executeUnit_jump_branch_info_branch_target = jump_branch_info_branch_target; // @[playground/src/pipeline/execute/ExecuteStage.scala 59:35]
  assign io_executeUnit_jump_branch_info_update_pht_index = jump_branch_info_update_pht_index; // @[playground/src/pipeline/execute/ExecuteStage.scala 59:35]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_pc <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_pc <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_pc <= io_decodeUnit_inst_0_pc; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_valid <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_valid <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_valid <= io_decodeUnit_inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_fusel <= 3'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_fusel <= 3'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_fusel <= io_decodeUnit_inst_0_info_fusel; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_op <= 7'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_op <= 7'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_op <= io_decodeUnit_inst_0_info_op; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_reg_wen <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_reg_wen <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_reg_wen <= io_decodeUnit_inst_0_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_reg_waddr <= io_decodeUnit_inst_0_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_imm <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_imm <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_imm <= io_decodeUnit_inst_0_info_imm; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_info_inst <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_info_inst <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_info_inst <= io_decodeUnit_inst_0_info_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_src_info_src1_data <= io_decodeUnit_inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_src_info_src2_data <= io_decodeUnit_inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_0 <= io_decodeUnit_inst_0_ex_exception_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_1 <= io_decodeUnit_inst_0_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_2 <= io_decodeUnit_inst_0_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_3 <= io_decodeUnit_inst_0_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_8 <= io_decodeUnit_inst_0_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_9 <= io_decodeUnit_inst_0_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_11 <= io_decodeUnit_inst_0_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_exception_12 <= io_decodeUnit_inst_0_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_0 <= io_decodeUnit_inst_0_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_1 <= io_decodeUnit_inst_0_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_2 <= io_decodeUnit_inst_0_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_3 <= io_decodeUnit_inst_0_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_4 <= io_decodeUnit_inst_0_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_5 <= io_decodeUnit_inst_0_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_6 <= io_decodeUnit_inst_0_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_7 <= io_decodeUnit_inst_0_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_8 <= io_decodeUnit_inst_0_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_9 <= io_decodeUnit_inst_0_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_10 <= io_decodeUnit_inst_0_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_interrupt_11 <= io_decodeUnit_inst_0_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_tval_0 <= io_decodeUnit_inst_0_ex_tval_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_tval_1 <= io_decodeUnit_inst_0_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_tval_2 <= io_decodeUnit_inst_0_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_0_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_0_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_0_ex_tval_12 <= io_decodeUnit_inst_0_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_pc <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_pc <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_pc <= io_decodeUnit_inst_1_pc; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_valid <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_valid <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_valid <= io_decodeUnit_inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_fusel <= 3'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_fusel <= 3'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_fusel <= io_decodeUnit_inst_1_info_fusel; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_op <= 7'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_op <= 7'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_op <= io_decodeUnit_inst_1_info_op; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_reg_wen <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_reg_wen <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_reg_wen <= io_decodeUnit_inst_1_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_reg_waddr <= io_decodeUnit_inst_1_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_imm <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_imm <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_imm <= io_decodeUnit_inst_1_info_imm; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_info_inst <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_info_inst <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_info_inst <= io_decodeUnit_inst_1_info_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_src_info_src1_data <= io_decodeUnit_inst_1_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_src_info_src2_data <= io_decodeUnit_inst_1_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_0 <= io_decodeUnit_inst_1_ex_exception_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_1 <= io_decodeUnit_inst_1_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_2 <= io_decodeUnit_inst_1_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_3 <= io_decodeUnit_inst_1_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_8 <= io_decodeUnit_inst_1_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_9 <= io_decodeUnit_inst_1_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_11 <= io_decodeUnit_inst_1_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_exception_12 <= io_decodeUnit_inst_1_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_0 <= io_decodeUnit_inst_1_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_1 <= io_decodeUnit_inst_1_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_2 <= io_decodeUnit_inst_1_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_3 <= io_decodeUnit_inst_1_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_4 <= io_decodeUnit_inst_1_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_5 <= io_decodeUnit_inst_1_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_6 <= io_decodeUnit_inst_1_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_7 <= io_decodeUnit_inst_1_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_8 <= io_decodeUnit_inst_1_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_9 <= io_decodeUnit_inst_1_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_10 <= io_decodeUnit_inst_1_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_interrupt_11 <= io_decodeUnit_inst_1_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_tval_0 <= io_decodeUnit_inst_1_ex_tval_0; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_tval_1 <= io_decodeUnit_inst_1_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_tval_2 <= io_decodeUnit_inst_1_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
      inst_1_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 40:63]
    end else if (io_ctrl_clear_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 44:28]
      inst_1_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 45:15]
    end else if (io_ctrl_allow_to_go_1) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 46:40]
      inst_1_ex_tval_12 <= io_decodeUnit_inst_1_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteStage.scala 47:15]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
      jump_branch_info_jump_regiser <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 52:26]
      jump_branch_info_jump_regiser <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 53:22]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 54:38]
      jump_branch_info_jump_regiser <= io_decodeUnit_jump_branch_info_jump_regiser; // @[playground/src/pipeline/execute/ExecuteStage.scala 55:22]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
      jump_branch_info_branch_inst <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 52:26]
      jump_branch_info_branch_inst <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 53:22]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 54:38]
      jump_branch_info_branch_inst <= io_decodeUnit_jump_branch_info_branch_inst; // @[playground/src/pipeline/execute/ExecuteStage.scala 55:22]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
      jump_branch_info_pred_branch <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 52:26]
      jump_branch_info_pred_branch <= 1'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 53:22]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 54:38]
      jump_branch_info_pred_branch <= io_decodeUnit_jump_branch_info_pred_branch; // @[playground/src/pipeline/execute/ExecuteStage.scala 55:22]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
      jump_branch_info_branch_target <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 52:26]
      jump_branch_info_branch_target <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 53:22]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 54:38]
      jump_branch_info_branch_target <= io_decodeUnit_jump_branch_info_branch_target; // @[playground/src/pipeline/execute/ExecuteStage.scala 55:22]
    end
    if (reset) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
      jump_branch_info_update_pht_index <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 41:33]
    end else if (io_ctrl_clear_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 52:26]
      jump_branch_info_update_pht_index <= 64'h0; // @[playground/src/pipeline/execute/ExecuteStage.scala 53:22]
    end else if (io_ctrl_allow_to_go_0) begin // @[playground/src/pipeline/execute/ExecuteStage.scala 54:38]
      jump_branch_info_update_pht_index <= io_decodeUnit_jump_branch_info_update_pht_index; // @[playground/src/pipeline/execute/ExecuteStage.scala 55:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  inst_0_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  inst_0_info_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_0_info_fusel = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  inst_0_info_op = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  inst_0_info_reg_wen = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  inst_0_info_reg_waddr = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  inst_0_info_imm = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  inst_0_info_inst = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  inst_0_src_info_src1_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  inst_0_src_info_src2_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  inst_0_ex_exception_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inst_0_ex_exception_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inst_0_ex_exception_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inst_0_ex_exception_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inst_0_ex_exception_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inst_0_ex_exception_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  inst_0_ex_exception_11 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  inst_0_ex_exception_12 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  inst_0_ex_interrupt_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  inst_0_ex_interrupt_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inst_0_ex_interrupt_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  inst_0_ex_interrupt_3 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  inst_0_ex_interrupt_4 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  inst_0_ex_interrupt_5 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  inst_0_ex_interrupt_6 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  inst_0_ex_interrupt_7 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  inst_0_ex_interrupt_8 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  inst_0_ex_interrupt_9 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  inst_0_ex_interrupt_10 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inst_0_ex_interrupt_11 = _RAND_29[0:0];
  _RAND_30 = {2{`RANDOM}};
  inst_0_ex_tval_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  inst_0_ex_tval_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  inst_0_ex_tval_2 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  inst_0_ex_tval_12 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  inst_1_pc = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  inst_1_info_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  inst_1_info_fusel = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  inst_1_info_op = _RAND_37[6:0];
  _RAND_38 = {1{`RANDOM}};
  inst_1_info_reg_wen = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  inst_1_info_reg_waddr = _RAND_39[4:0];
  _RAND_40 = {2{`RANDOM}};
  inst_1_info_imm = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  inst_1_info_inst = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  inst_1_src_info_src1_data = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  inst_1_src_info_src2_data = _RAND_43[63:0];
  _RAND_44 = {1{`RANDOM}};
  inst_1_ex_exception_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  inst_1_ex_exception_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  inst_1_ex_exception_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  inst_1_ex_exception_3 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  inst_1_ex_exception_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  inst_1_ex_exception_9 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  inst_1_ex_exception_11 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  inst_1_ex_exception_12 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  inst_1_ex_interrupt_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  inst_1_ex_interrupt_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  inst_1_ex_interrupt_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  inst_1_ex_interrupt_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  inst_1_ex_interrupt_4 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  inst_1_ex_interrupt_5 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  inst_1_ex_interrupt_6 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  inst_1_ex_interrupt_7 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  inst_1_ex_interrupt_8 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  inst_1_ex_interrupt_9 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  inst_1_ex_interrupt_10 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  inst_1_ex_interrupt_11 = _RAND_63[0:0];
  _RAND_64 = {2{`RANDOM}};
  inst_1_ex_tval_0 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  inst_1_ex_tval_1 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  inst_1_ex_tval_2 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  inst_1_ex_tval_12 = _RAND_67[63:0];
  _RAND_68 = {1{`RANDOM}};
  jump_branch_info_jump_regiser = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  jump_branch_info_branch_inst = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  jump_branch_info_pred_branch = _RAND_70[0:0];
  _RAND_71 = {2{`RANDOM}};
  jump_branch_info_branch_target = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  jump_branch_info_update_pht_index = _RAND_72[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Alu(
  input  [6:0]  io_info_op, // @[playground/src/pipeline/execute/fu/Alu.scala 9:14]
  input  [63:0] io_src_info_src1_data, // @[playground/src/pipeline/execute/fu/Alu.scala 9:14]
  input  [63:0] io_src_info_src2_data, // @[playground/src/pipeline/execute/fu/Alu.scala 9:14]
  output [63:0] io_result // @[playground/src/pipeline/execute/fu/Alu.scala 9:14]
);
  wire  is_sub = ~io_info_op[5]; // @[playground/src/pipeline/execute/fu/Alu.scala 17:16]
  wire [63:0] _sum_T_1 = is_sub ? 64'hffffffffffffffff : 64'h0; // @[playground/src/pipeline/execute/fu/Alu.scala 18:37]
  wire [63:0] _sum_T_2 = io_src_info_src2_data ^ _sum_T_1; // @[playground/src/pipeline/execute/fu/Alu.scala 18:31]
  wire [64:0] _sum_T_3 = io_src_info_src1_data + _sum_T_2; // @[playground/src/pipeline/execute/fu/Alu.scala 18:22]
  wire [64:0] _GEN_0 = {{64'd0}, is_sub}; // @[playground/src/pipeline/execute/fu/Alu.scala 18:54]
  wire [64:0] sum = _sum_T_3 + _GEN_0; // @[playground/src/pipeline/execute/fu/Alu.scala 18:54]
  wire [63:0] xor_ = io_src_info_src1_data ^ io_src_info_src2_data; // @[playground/src/pipeline/execute/fu/Alu.scala 19:21]
  wire  sltu = ~sum[64]; // @[playground/src/pipeline/execute/fu/Alu.scala 20:16]
  wire  slt = xor_[63] ^ sltu; // @[playground/src/pipeline/execute/fu/Alu.scala 21:30]
  wire [63:0] _shsrc1_T_2 = {32'h0,io_src_info_src1_data[31:0]}; // @[playground/src/defines/Util.scala 41:44]
  wire  shsrc1_signBit = io_src_info_src1_data[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _shsrc1_T_5 = shsrc1_signBit ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _shsrc1_T_6 = {_shsrc1_T_5,io_src_info_src1_data[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire [63:0] _shsrc1_T_8 = 7'h15 == io_info_op ? _shsrc1_T_2 : io_src_info_src1_data; // @[playground/src/pipeline/execute/fu/Alu.scala 23:48]
  wire [63:0] shsrc1 = 7'h1d == io_info_op ? _shsrc1_T_6 : _shsrc1_T_8; // @[playground/src/pipeline/execute/fu/Alu.scala 23:48]
  wire [5:0] shamt = io_info_op[4] ? {{1'd0}, io_src_info_src2_data[4:0]} : io_src_info_src2_data[5:0]; // @[playground/src/pipeline/execute/fu/Alu.scala 29:18]
  wire [126:0] _GEN_1 = {{63'd0}, shsrc1}; // @[playground/src/pipeline/execute/fu/Alu.scala 32:34]
  wire [126:0] _res_T_1 = _GEN_1 << shamt; // @[playground/src/pipeline/execute/fu/Alu.scala 32:34]
  wire [63:0] _res_T_3 = {63'h0,slt}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _res_T_4 = {63'h0,sltu}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _res_T_5 = shsrc1 >> shamt; // @[playground/src/pipeline/execute/fu/Alu.scala 36:33]
  wire [63:0] _res_T_6 = io_src_info_src1_data | io_src_info_src2_data; // @[playground/src/pipeline/execute/fu/Alu.scala 37:31]
  wire [63:0] _res_T_7 = io_src_info_src1_data & io_src_info_src2_data; // @[playground/src/pipeline/execute/fu/Alu.scala 38:31]
  wire [63:0] _res_T_8 = 7'h1d == io_info_op ? _shsrc1_T_6 : _shsrc1_T_8; // @[playground/src/pipeline/execute/fu/Alu.scala 39:34]
  wire [63:0] _res_T_10 = $signed(_res_T_8) >>> shamt; // @[playground/src/pipeline/execute/fu/Alu.scala 39:51]
  wire [64:0] _res_T_12 = 4'h1 == io_info_op[3:0] ? {{1'd0}, _res_T_1[63:0]} : sum; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] _res_T_14 = 4'h2 == io_info_op[3:0] ? {{1'd0}, _res_T_3} : _res_T_12; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] _res_T_16 = 4'h3 == io_info_op[3:0] ? {{1'd0}, _res_T_4} : _res_T_14; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] _res_T_18 = 4'h4 == io_info_op[3:0] ? {{1'd0}, xor_} : _res_T_16; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] _res_T_20 = 4'h5 == io_info_op[3:0] ? {{1'd0}, _res_T_5} : _res_T_18; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] _res_T_22 = 4'h6 == io_info_op[3:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] _res_T_24 = 4'h7 == io_info_op[3:0] ? {{1'd0}, _res_T_7} : _res_T_22; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire [64:0] res = 4'hd == io_info_op[3:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[playground/src/pipeline/execute/fu/Alu.scala 30:37]
  wire  io_result_signBit = res[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _io_result_T_3 = io_result_signBit ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_result_T_4 = {_io_result_T_3,res[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire [64:0] _io_result_T_5 = io_info_op[4] ? {{1'd0}, _io_result_T_4} : res; // @[playground/src/pipeline/execute/fu/Alu.scala 42:19]
  assign io_result = _io_result_T_5[63:0]; // @[playground/src/pipeline/execute/fu/Alu.scala 42:13]
endmodule
module BranchCtrl(
  input  [63:0] io_in_pc, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input         io_in_info_valid, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input  [2:0]  io_in_info_fusel, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input  [6:0]  io_in_info_op, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input  [63:0] io_in_src_info_src1_data, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input  [63:0] io_in_src_info_src2_data, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input         io_in_pred_branch, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input         io_in_jump_regiser, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  input  [63:0] io_in_branch_target, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  output        io_out_branch, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  output        io_out_pred_fail, // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
  output [63:0] io_out_target // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 9:14]
);
  wire  _valid_T_2 = ~io_in_info_op[3]; // @[playground/src/defines/isa/Instructions.scala 74:36]
  wire  valid = io_in_info_fusel == 3'h5 & _valid_T_2 & io_in_info_valid; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 25:74]
  wire  _is_sub_T_2 = ~_valid_T_2; // @[playground/src/defines/isa/Instructions.scala 75:36]
  wire  is_sub = ~_is_sub_T_2; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 29:16]
  wire [63:0] _adder_T_1 = is_sub ? 64'hffffffffffffffff : 64'h0; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 30:37]
  wire [63:0] _adder_T_2 = io_in_src_info_src2_data ^ _adder_T_1; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 30:31]
  wire [64:0] _adder_T_3 = io_in_src_info_src1_data + _adder_T_2; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 30:22]
  wire [64:0] _GEN_0 = {{64'd0}, is_sub}; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 30:54]
  wire [64:0] adder = _adder_T_3 + _GEN_0; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 30:54]
  wire [63:0] xor_ = io_in_src_info_src1_data ^ io_in_src_info_src2_data; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 31:21]
  wire  sltu = ~adder[64]; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 32:16]
  wire  slt = xor_[63] ^ sltu; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 33:30]
  wire  _T_1 = ~(|xor_); // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 35:48]
  wire  _io_out_branch_T_1 = 2'h0 == io_in_info_op[2:1]; // @[playground/src/defines/Util.scala 46:34]
  wire  _io_out_branch_T_2 = 2'h2 == io_in_info_op[2:1]; // @[playground/src/defines/Util.scala 46:34]
  wire  _io_out_branch_T_3 = 2'h3 == io_in_info_op[2:1]; // @[playground/src/defines/Util.scala 46:34]
  wire  _io_out_branch_T_8 = _io_out_branch_T_1 & _T_1 | _io_out_branch_T_2 & slt | _io_out_branch_T_3 & sltu; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_out_target_T = io_out_pred_fail & io_out_branch; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 44:25]
  wire  _io_out_target_T_2 = io_out_pred_fail & ~io_out_branch; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 45:25]
  wire [63:0] _io_out_target_T_4 = io_in_pc + 64'h4; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 45:57]
  wire [63:0] _io_out_target_T_6 = io_in_src_info_src1_data + io_in_src_info_src2_data; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 46:54]
  wire [63:0] _io_out_target_T_8 = _io_out_target_T_6 & 64'hfffffffffffffffe; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 46:62]
  wire [63:0] _io_out_target_T_9 = _io_out_target_T ? io_in_branch_target : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_target_T_10 = _io_out_target_T_2 ? _io_out_target_T_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_target_T_11 = io_in_jump_regiser ? _io_out_target_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_target_T_12 = _io_out_target_T_9 | _io_out_target_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_branch = (_io_out_branch_T_8 ^ io_in_info_op[0]) & valid; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 41:85]
  assign io_out_pred_fail = io_in_pred_branch != io_out_branch; // @[playground/src/pipeline/execute/fu/BranchCtrl.scala 39:41]
  assign io_out_target = _io_out_target_T_12 | _io_out_target_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
endmodule
module Mul(
  input          clock,
  input          reset,
  input  [64:0]  io_src1, // @[playground/src/pipeline/execute/fu/Mul.scala 21:14]
  input  [64:0]  io_src2, // @[playground/src/pipeline/execute/fu/Mul.scala 21:14]
  input          io_en, // @[playground/src/pipeline/execute/fu/Mul.scala 21:14]
  input          io_allow_to_go, // @[playground/src/pipeline/execute/fu/Mul.scala 21:14]
  output         io_ready, // @[playground/src/pipeline/execute/fu/Mul.scala 21:14]
  output [127:0] io_result // @[playground/src/pipeline/execute/fu/Mul.scala 21:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] cnt; // @[playground/src/pipeline/execute/fu/Mul.scala 52:22]
  wire  _cnt_T_1 = io_en & ~io_ready; // @[playground/src/pipeline/execute/fu/Mul.scala 56:16]
  wire [1:0] _cnt_T_3 = cnt + 2'h1; // @[playground/src/pipeline/execute/fu/Mul.scala 56:38]
  reg [127:0] signed_; // @[playground/src/pipeline/execute/fu/Mul.scala 61:25]
  wire [129:0] _signed_T_3 = $signed(io_src1) * $signed(io_src2); // @[playground/src/pipeline/execute/fu/Mul.scala 63:51]
  wire [129:0] _GEN_0 = io_en ? _signed_T_3 : {{2'd0}, signed_}; // @[playground/src/pipeline/execute/fu/Mul.scala 62:17 63:14 61:25]
  wire [129:0] _GEN_1 = reset ? 130'h0 : _GEN_0; // @[playground/src/pipeline/execute/fu/Mul.scala 61:{25,25}]
  assign io_ready = cnt >= 2'h2; // @[playground/src/pipeline/execute/fu/Mul.scala 66:22]
  assign io_result = signed_; // @[playground/src/pipeline/execute/fu/Mul.scala 65:15]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/execute/fu/Mul.scala 52:22]
      cnt <= 2'h0; // @[playground/src/pipeline/execute/fu/Mul.scala 52:22]
    end else if (_cnt_T_1) begin // @[src/main/scala/chisel3/util/Mux.scala 141:16]
      cnt <= _cnt_T_3;
    end else if (io_allow_to_go) begin // @[src/main/scala/chisel3/util/Mux.scala 141:16]
      cnt <= 2'h0;
    end
    signed_ <= _GEN_1[127:0]; // @[playground/src/pipeline/execute/fu/Mul.scala 61:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[1:0];
  _RAND_1 = {4{`RANDOM}};
  signed_ = _RAND_1[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Div(
  input          clock,
  input          reset,
  input  [63:0]  io_src1, // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
  input  [63:0]  io_src2, // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
  input          io_signed, // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
  input          io_en, // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
  input          io_allow_to_go, // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
  output         io_ready, // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
  output [127:0] io_result // @[playground/src/pipeline/execute/fu/Div.scala 44:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] cnt; // @[playground/src/pipeline/execute/fu/Div.scala 127:22]
  wire  _cnt_T_1 = io_en & ~io_ready; // @[playground/src/pipeline/execute/fu/Div.scala 131:16]
  wire [3:0] _cnt_T_3 = cnt + 4'h1; // @[playground/src/pipeline/execute/fu/Div.scala 131:38]
  wire  dividend_signed = io_src1[63] & io_signed; // @[playground/src/pipeline/execute/fu/Div.scala 138:45]
  wire  divisor_signed = io_src2[63] & io_signed; // @[playground/src/pipeline/execute/fu/Div.scala 139:45]
  wire [63:0] _dividend_abs_T_1 = 64'h0 - io_src1; // @[playground/src/pipeline/execute/fu/Div.scala 141:46]
  wire [63:0] dividend_abs = dividend_signed ? _dividend_abs_T_1 : io_src1; // @[playground/src/pipeline/execute/fu/Div.scala 141:27]
  wire [63:0] _divisor_abs_T_1 = 64'h0 - io_src2; // @[playground/src/pipeline/execute/fu/Div.scala 142:45]
  wire [63:0] divisor_abs = divisor_signed ? _divisor_abs_T_1 : io_src2; // @[playground/src/pipeline/execute/fu/Div.scala 142:27]
  wire  quotient_signed = (io_src1[63] ^ io_src2[63]) & io_signed; // @[playground/src/pipeline/execute/fu/Div.scala 144:68]
  wire [63:0] quotient_abs = dividend_abs / divisor_abs; // @[playground/src/pipeline/execute/fu/Div.scala 147:38]
  wire [127:0] _remainder_abs_T = quotient_abs * divisor_abs; // @[playground/src/pipeline/execute/fu/Div.scala 148:53]
  wire [127:0] _GEN_4 = {{64'd0}, dividend_abs}; // @[playground/src/pipeline/execute/fu/Div.scala 148:38]
  wire [127:0] remainder_abs = _GEN_4 - _remainder_abs_T; // @[playground/src/pipeline/execute/fu/Div.scala 148:38]
  reg [63:0] quotient; // @[playground/src/pipeline/execute/fu/Div.scala 150:28]
  reg [63:0] remainder; // @[playground/src/pipeline/execute/fu/Div.scala 151:28]
  wire [63:0] _quotient_T_2 = 64'h0 - quotient_abs; // @[playground/src/pipeline/execute/fu/Div.scala 154:57]
  wire [63:0] _quotient_T_3 = dividend_abs / divisor_abs; // @[playground/src/pipeline/execute/fu/Div.scala 154:78]
  wire [127:0] _remainder_T_2 = 128'h0 - remainder_abs; // @[playground/src/pipeline/execute/fu/Div.scala 155:59]
  wire [127:0] _remainder_T_3 = _GEN_4 - _remainder_abs_T; // @[playground/src/pipeline/execute/fu/Div.scala 155:81]
  wire [127:0] _remainder_T_4 = dividend_signed ? $signed(_remainder_T_2) : $signed(_remainder_T_3); // @[playground/src/pipeline/execute/fu/Div.scala 155:23]
  wire [63:0] _remainder_T_5 = io_src1; // @[playground/src/pipeline/execute/fu/Div.scala 158:30]
  wire [127:0] _GEN_1 = io_src2 == 64'h0 ? $signed({{64{_remainder_T_5[63]}},_remainder_T_5}) : $signed(_remainder_T_4); // @[playground/src/pipeline/execute/fu/Div.scala 155:17 156:29 158:19]
  wire [127:0] _GEN_3 = io_en ? $signed(_GEN_1) : $signed({{64{remainder[63]}},remainder}); // @[playground/src/pipeline/execute/fu/Div.scala 153:17 151:28]
  wire [127:0] _GEN_5 = reset ? $signed(128'sh0) : $signed(_GEN_3); // @[playground/src/pipeline/execute/fu/Div.scala 151:{28,28}]
  assign io_ready = cnt >= 4'h8; // @[playground/src/pipeline/execute/fu/Div.scala 162:22]
  assign io_result = {remainder,quotient}; // @[playground/src/pipeline/execute/fu/Div.scala 163:21]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/execute/fu/Div.scala 127:22]
      cnt <= 4'h0; // @[playground/src/pipeline/execute/fu/Div.scala 127:22]
    end else if (_cnt_T_1) begin // @[src/main/scala/chisel3/util/Mux.scala 141:16]
      cnt <= _cnt_T_3;
    end else if (io_allow_to_go) begin // @[src/main/scala/chisel3/util/Mux.scala 141:16]
      cnt <= 4'h0;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Div.scala 150:28]
      quotient <= 64'sh0; // @[playground/src/pipeline/execute/fu/Div.scala 150:28]
    end else if (io_en) begin // @[playground/src/pipeline/execute/fu/Div.scala 153:17]
      if (io_src2 == 64'h0) begin // @[playground/src/pipeline/execute/fu/Div.scala 156:29]
        quotient <= -64'sh1; // @[playground/src/pipeline/execute/fu/Div.scala 157:19]
      end else if (quotient_signed) begin // @[playground/src/pipeline/execute/fu/Div.scala 154:23]
        quotient <= _quotient_T_2;
      end else begin
        quotient <= _quotient_T_3;
      end
    end
    remainder <= _GEN_5[63:0]; // @[playground/src/pipeline/execute/fu/Div.scala 151:{28,28}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[3:0];
  _RAND_1 = {2{`RANDOM}};
  quotient = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  remainder = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mdu(
  input         clock,
  input         reset,
  input         io_info_valid, // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
  input  [6:0]  io_info_op, // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
  input  [63:0] io_src_info_src1_data, // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
  input  [63:0] io_src_info_src2_data, // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
  input         io_allow_to_go, // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
  output        io_ready, // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
  output [63:0] io_result // @[playground/src/pipeline/execute/fu/Mdu.scala 10:14]
);
  wire  Mul_clock; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire  Mul_reset; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire [64:0] Mul_io_src1; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire [64:0] Mul_io_src2; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire  Mul_io_en; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire  Mul_io_allow_to_go; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire  Mul_io_ready; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire [127:0] Mul_io_result; // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
  wire  Div_clock; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire  Div_reset; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire [63:0] Div_io_src1; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire [63:0] Div_io_src2; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire  Div_io_signed; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire  Div_io_en; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire  Div_io_allow_to_go; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire  Div_io_ready; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire [127:0] Div_io_result; // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
  wire  is_div = io_info_op[2]; // @[playground/src/defines/isa/Instructions.scala 140:31]
  wire  is_w = io_info_op[3]; // @[playground/src/defines/isa/Instructions.scala 142:31]
  wire [64:0] _T_1 = {1'h0,io_src_info_src1_data}; // @[playground/src/defines/Util.scala 41:44]
  wire  signBit = io_src_info_src1_data[63]; // @[playground/src/defines/Util.scala 33:20]
  wire [64:0] _T_2 = {signBit,io_src_info_src1_data}; // @[playground/src/defines/Util.scala 34:44]
  wire  _T_5 = 2'h0 == io_info_op[1:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _T_6 = 2'h1 == io_info_op[1:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _T_7 = 2'h2 == io_info_op[1:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _T_8 = 2'h3 == io_info_op[1:0]; // @[playground/src/defines/Util.scala 46:34]
  wire [64:0] _T_9 = _T_5 ? _T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_10 = _T_6 ? _T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_11 = _T_7 ? _T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_12 = _T_8 ? _T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_13 = _T_9 | _T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_14 = _T_13 | _T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_17 = {1'h0,io_src_info_src2_data}; // @[playground/src/defines/Util.scala 41:44]
  wire  signBit_2 = io_src_info_src2_data[63]; // @[playground/src/defines/Util.scala 33:20]
  wire [64:0] _T_18 = {signBit_2,io_src_info_src2_data}; // @[playground/src/defines/Util.scala 34:44]
  wire [64:0] _T_25 = _T_5 ? _T_17 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_26 = _T_6 ? _T_18 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_27 = _T_7 ? _T_17 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_28 = _T_8 ? _T_17 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_29 = _T_25 | _T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _T_30 = _T_29 | _T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_37 = is_div & ~io_info_op[0]; // @[playground/src/defines/isa/Instructions.scala 141:39]
  wire  signBit_3 = io_src_info_src1_data[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _T_40 = signBit_3 ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _T_41 = {_T_40,io_src_info_src1_data[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire [63:0] _T_43 = {32'h0,io_src_info_src1_data[31:0]}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _T_44 = _T_37 ? _T_41 : _T_43; // @[playground/src/pipeline/execute/fu/Mdu.scala 45:18]
  wire  signBit_4 = io_src_info_src2_data[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _T_52 = signBit_4 ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _T_53 = {_T_52,io_src_info_src2_data[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire [63:0] _T_55 = {32'h0,io_src_info_src2_data[31:0]}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _T_56 = _T_37 ? _T_53 : _T_55; // @[playground/src/pipeline/execute/fu/Mdu.scala 45:18]
  wire [63:0] mul_result = io_info_op[1:0] == 2'h0 ? Mul_io_result[63:0] : Mul_io_result[127:64]; // @[playground/src/pipeline/execute/fu/Mdu.scala 52:23]
  wire [63:0] div_result = io_info_op[1] ? Div_io_result[127:64] : Div_io_result[63:0]; // @[playground/src/pipeline/execute/fu/Mdu.scala 53:23]
  wire [63:0] result = is_div ? div_result : mul_result; // @[playground/src/pipeline/execute/fu/Mdu.scala 54:23]
  wire  io_result_signBit = result[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _io_result_T_2 = io_result_signBit ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_result_T_3 = {_io_result_T_2,result[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  Mul Mul ( // @[playground/src/pipeline/execute/fu/Mdu.scala 19:19]
    .clock(Mul_clock),
    .reset(Mul_reset),
    .io_src1(Mul_io_src1),
    .io_src2(Mul_io_src2),
    .io_en(Mul_io_en),
    .io_allow_to_go(Mul_io_allow_to_go),
    .io_ready(Mul_io_ready),
    .io_result(Mul_io_result)
  );
  Div Div ( // @[playground/src/pipeline/execute/fu/Mdu.scala 20:19]
    .clock(Div_clock),
    .reset(Div_reset),
    .io_src1(Div_io_src1),
    .io_src2(Div_io_src2),
    .io_signed(Div_io_signed),
    .io_en(Div_io_en),
    .io_allow_to_go(Div_io_allow_to_go),
    .io_ready(Div_io_ready),
    .io_result(Div_io_result)
  );
  assign io_ready = is_div ? Div_io_ready : Mul_io_ready; // @[playground/src/pipeline/execute/fu/Mdu.scala 56:19]
  assign io_result = is_w ? _io_result_T_3 : result; // @[playground/src/pipeline/execute/fu/Mdu.scala 57:19]
  assign Mul_clock = clock;
  assign Mul_reset = reset;
  assign Mul_io_src1 = _T_14 | _T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Mul_io_src2 = _T_30 | _T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Mul_io_en = io_info_valid & ~is_div; // @[playground/src/pipeline/execute/fu/Mdu.scala 41:28]
  assign Mul_io_allow_to_go = io_allow_to_go; // @[playground/src/pipeline/execute/fu/Mdu.scala 42:19]
  assign Div_clock = clock;
  assign Div_reset = reset;
  assign Div_io_src1 = is_w ? _T_44 : io_src_info_src1_data; // @[playground/src/pipeline/execute/fu/Mdu.scala 45:8]
  assign Div_io_src2 = is_w ? _T_56 : io_src_info_src2_data; // @[playground/src/pipeline/execute/fu/Mdu.scala 45:8]
  assign Div_io_signed = is_div & ~io_info_op[0]; // @[playground/src/defines/isa/Instructions.scala 141:39]
  assign Div_io_en = io_info_valid & is_div; // @[playground/src/pipeline/execute/fu/Mdu.scala 49:28]
  assign Div_io_allow_to_go = io_allow_to_go; // @[playground/src/pipeline/execute/fu/Mdu.scala 50:19]
endmodule
module Fu(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output        io_ctrl_stall, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_0_pc, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input         io_inst_0_info_valid, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [2:0]  io_inst_0_info_fusel, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [6:0]  io_inst_0_info_op, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_0_info_imm, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_0_src_info_src1_data, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_0_src_info_src2_data, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output [63:0] io_inst_0_result_mdu, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output [63:0] io_inst_0_result_alu, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input         io_inst_1_info_valid, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [2:0]  io_inst_1_info_fusel, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [6:0]  io_inst_1_info_op, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_1_info_imm, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_1_src_info_src1_data, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_inst_1_src_info_src2_data, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output [63:0] io_inst_1_result_mdu, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output [63:0] io_inst_1_result_alu, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output [63:0] io_dataMemory_addr, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input         io_branch_pred_branch, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input         io_branch_jump_regiser, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  input  [63:0] io_branch_branch_target, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output        io_branch_branch, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output        io_branch_flush, // @[playground/src/pipeline/execute/Fu.scala 10:14]
  output [63:0] io_branch_target // @[playground/src/pipeline/execute/Fu.scala 10:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] alu_0_io_info_op; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] alu_0_io_src_info_src1_data; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] alu_0_io_src_info_src2_data; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] alu_0_io_result; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [6:0] alu_1_io_info_op; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] alu_1_io_src_info_src1_data; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] alu_1_io_src_info_src2_data; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] alu_1_io_result; // @[playground/src/pipeline/execute/Fu.scala 37:57]
  wire [63:0] BranchCtrl_io_in_pc; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire  BranchCtrl_io_in_info_valid; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire [2:0] BranchCtrl_io_in_info_fusel; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire [6:0] BranchCtrl_io_in_info_op; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire [63:0] BranchCtrl_io_in_src_info_src1_data; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire [63:0] BranchCtrl_io_in_src_info_src2_data; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire  BranchCtrl_io_in_pred_branch; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire  BranchCtrl_io_in_jump_regiser; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire [63:0] BranchCtrl_io_in_branch_target; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire  BranchCtrl_io_out_branch; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire  BranchCtrl_io_out_pred_fail; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire [63:0] BranchCtrl_io_out_target; // @[playground/src/pipeline/execute/Fu.scala 38:26]
  wire  Mdu_clock; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire  Mdu_reset; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire  Mdu_io_info_valid; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire [6:0] Mdu_io_info_op; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire [63:0] Mdu_io_src_info_src1_data; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire [63:0] Mdu_io_src_info_src2_data; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire  Mdu_io_allow_to_go; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire  Mdu_io_ready; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire [63:0] Mdu_io_result; // @[playground/src/pipeline/execute/Fu.scala 39:26]
  wire  _alu_0_io_info_T = io_inst_0_info_fusel == 3'h0; // @[playground/src/pipeline/execute/Fu.scala 54:53]
  wire  _alu_1_io_info_T = io_inst_1_info_fusel == 3'h0; // @[playground/src/pipeline/execute/Fu.scala 54:53]
  wire  mdu_sel_0 = io_inst_0_info_fusel == 3'h2; // @[playground/src/pipeline/execute/Fu.scala 59:27]
  wire  mdu_sel_1 = io_inst_1_info_fusel == 3'h2; // @[playground/src/pipeline/execute/Fu.scala 60:27]
  wire [6:0] _T_op = mdu_sel_1 ? io_inst_1_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _T_2_src1_data = mdu_sel_1 ? io_inst_1_src_info_src1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _T_2_src2_data = mdu_sel_1 ? io_inst_1_src_info_src2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _mem_addr_T_2 = io_inst_0_src_info_src1_data + io_inst_0_info_imm; // @[playground/src/pipeline/execute/Fu.scala 85:37]
  wire [63:0] mem_addr_0 = io_inst_0_info_op[5] ? io_inst_0_src_info_src1_data : _mem_addr_T_2; // @[playground/src/pipeline/execute/Fu.scala 82:8]
  wire [63:0] _mem_addr_T_5 = io_inst_1_src_info_src1_data + io_inst_1_info_imm; // @[playground/src/pipeline/execute/Fu.scala 85:37]
  wire [63:0] mem_addr_1 = io_inst_1_info_op[5] ? io_inst_1_src_info_src1_data : _mem_addr_T_5; // @[playground/src/pipeline/execute/Fu.scala 82:8]
  reg [63:0] mem_addr_last; // @[playground/src/pipeline/execute/Fu.scala 89:32]
  wire  _io_dataMemory_addr_T = ~io_ctrl_allow_to_go; // @[playground/src/pipeline/execute/Fu.scala 91:5]
  wire [63:0] _io_dataMemory_addr_T_2 = io_inst_0_info_fusel == 3'h1 ? mem_addr_0 : mem_addr_1; // @[playground/src/pipeline/execute/Fu.scala 93:8]
  Alu alu_0 ( // @[playground/src/pipeline/execute/Fu.scala 37:57]
    .io_info_op(alu_0_io_info_op),
    .io_src_info_src1_data(alu_0_io_src_info_src1_data),
    .io_src_info_src2_data(alu_0_io_src_info_src2_data),
    .io_result(alu_0_io_result)
  );
  Alu alu_1 ( // @[playground/src/pipeline/execute/Fu.scala 37:57]
    .io_info_op(alu_1_io_info_op),
    .io_src_info_src1_data(alu_1_io_src_info_src1_data),
    .io_src_info_src2_data(alu_1_io_src_info_src2_data),
    .io_result(alu_1_io_result)
  );
  BranchCtrl BranchCtrl ( // @[playground/src/pipeline/execute/Fu.scala 38:26]
    .io_in_pc(BranchCtrl_io_in_pc),
    .io_in_info_valid(BranchCtrl_io_in_info_valid),
    .io_in_info_fusel(BranchCtrl_io_in_info_fusel),
    .io_in_info_op(BranchCtrl_io_in_info_op),
    .io_in_src_info_src1_data(BranchCtrl_io_in_src_info_src1_data),
    .io_in_src_info_src2_data(BranchCtrl_io_in_src_info_src2_data),
    .io_in_pred_branch(BranchCtrl_io_in_pred_branch),
    .io_in_jump_regiser(BranchCtrl_io_in_jump_regiser),
    .io_in_branch_target(BranchCtrl_io_in_branch_target),
    .io_out_branch(BranchCtrl_io_out_branch),
    .io_out_pred_fail(BranchCtrl_io_out_pred_fail),
    .io_out_target(BranchCtrl_io_out_target)
  );
  Mdu Mdu ( // @[playground/src/pipeline/execute/Fu.scala 39:26]
    .clock(Mdu_clock),
    .reset(Mdu_reset),
    .io_info_valid(Mdu_io_info_valid),
    .io_info_op(Mdu_io_info_op),
    .io_src_info_src1_data(Mdu_io_src_info_src1_data),
    .io_src_info_src2_data(Mdu_io_src_info_src2_data),
    .io_allow_to_go(Mdu_io_allow_to_go),
    .io_ready(Mdu_io_ready),
    .io_result(Mdu_io_result)
  );
  assign io_ctrl_stall = (mdu_sel_0 | mdu_sel_1) & ~Mdu_io_ready; // @[playground/src/pipeline/execute/Fu.scala 73:76]
  assign io_inst_0_result_mdu = Mdu_io_result; // @[playground/src/pipeline/execute/Fu.scala 76:25]
  assign io_inst_0_result_alu = alu_0_io_result; // @[playground/src/pipeline/execute/Fu.scala 75:25]
  assign io_inst_1_result_mdu = Mdu_io_result; // @[playground/src/pipeline/execute/Fu.scala 79:25]
  assign io_inst_1_result_alu = alu_1_io_result; // @[playground/src/pipeline/execute/Fu.scala 78:25]
  assign io_dataMemory_addr = _io_dataMemory_addr_T ? mem_addr_last : _io_dataMemory_addr_T_2; // @[playground/src/pipeline/execute/Fu.scala 90:28]
  assign io_branch_branch = BranchCtrl_io_out_branch; // @[playground/src/pipeline/execute/Fu.scala 47:31]
  assign io_branch_flush = BranchCtrl_io_out_pred_fail | io_branch_jump_regiser; // @[playground/src/pipeline/execute/Fu.scala 49:52]
  assign io_branch_target = BranchCtrl_io_out_target; // @[playground/src/pipeline/execute/Fu.scala 51:20]
  assign alu_0_io_info_op = io_inst_0_info_fusel == 3'h0 ? io_inst_0_info_op : 7'h0; // @[playground/src/pipeline/execute/Fu.scala 54:30]
  assign alu_0_io_src_info_src1_data = _alu_0_io_info_T ? io_inst_0_src_info_src1_data : 64'h0; // @[playground/src/pipeline/execute/Fu.scala 55:30]
  assign alu_0_io_src_info_src2_data = _alu_0_io_info_T ? io_inst_0_src_info_src2_data : 64'h0; // @[playground/src/pipeline/execute/Fu.scala 55:30]
  assign alu_1_io_info_op = io_inst_1_info_fusel == 3'h0 ? io_inst_1_info_op : 7'h0; // @[playground/src/pipeline/execute/Fu.scala 54:30]
  assign alu_1_io_src_info_src1_data = _alu_1_io_info_T ? io_inst_1_src_info_src1_data : 64'h0; // @[playground/src/pipeline/execute/Fu.scala 55:30]
  assign alu_1_io_src_info_src2_data = _alu_1_io_info_T ? io_inst_1_src_info_src2_data : 64'h0; // @[playground/src/pipeline/execute/Fu.scala 55:30]
  assign BranchCtrl_io_in_pc = io_inst_0_pc; // @[playground/src/pipeline/execute/Fu.scala 41:31]
  assign BranchCtrl_io_in_info_valid = io_inst_0_info_valid; // @[playground/src/pipeline/execute/Fu.scala 42:31]
  assign BranchCtrl_io_in_info_fusel = io_inst_0_info_fusel; // @[playground/src/pipeline/execute/Fu.scala 42:31]
  assign BranchCtrl_io_in_info_op = io_inst_0_info_op; // @[playground/src/pipeline/execute/Fu.scala 42:31]
  assign BranchCtrl_io_in_src_info_src1_data = io_inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/Fu.scala 43:31]
  assign BranchCtrl_io_in_src_info_src2_data = io_inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/Fu.scala 43:31]
  assign BranchCtrl_io_in_pred_branch = io_branch_pred_branch; // @[playground/src/pipeline/execute/Fu.scala 44:31]
  assign BranchCtrl_io_in_jump_regiser = io_branch_jump_regiser; // @[playground/src/pipeline/execute/Fu.scala 45:31]
  assign BranchCtrl_io_in_branch_target = io_branch_branch_target; // @[playground/src/pipeline/execute/Fu.scala 46:31]
  assign Mdu_clock = clock;
  assign Mdu_reset = reset;
  assign Mdu_io_info_valid = mdu_sel_0 ? io_inst_0_info_valid : mdu_sel_1 & io_inst_1_info_valid; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign Mdu_io_info_op = mdu_sel_0 ? io_inst_0_info_op : _T_op; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign Mdu_io_src_info_src1_data = mdu_sel_0 ? io_inst_0_src_info_src1_data : _T_2_src1_data; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign Mdu_io_src_info_src2_data = mdu_sel_0 ? io_inst_0_src_info_src2_data : _T_2_src2_data; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign Mdu_io_allow_to_go = io_ctrl_allow_to_go; // @[playground/src/pipeline/execute/Fu.scala 71:19]
  always @(posedge clock) begin
    if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/execute/Fu.scala 89:32]
      mem_addr_last <= io_dataMemory_addr; // @[playground/src/pipeline/execute/Fu.scala 89:32]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mem_addr_last = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ExecuteUnit(
  input         clock,
  input         reset,
  output        io_ctrl_inst_0_is_load, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [4:0]  io_ctrl_inst_0_reg_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_ctrl_inst_1_is_load, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [4:0]  io_ctrl_inst_1_reg_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_ctrl_flush, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_ctrl_allow_to_go, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_ctrl_fu_allow_to_go, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_ctrl_fu_stall, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_pc, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_info_valid, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [2:0]  io_executeStage_inst_0_info_fusel, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [6:0]  io_executeStage_inst_0_info_op, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [4:0]  io_executeStage_inst_0_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_info_imm, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_info_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_0_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_0_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_pc, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_info_valid, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [2:0]  io_executeStage_inst_1_info_fusel, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [6:0]  io_executeStage_inst_1_info_op, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [4:0]  io_executeStage_inst_1_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_info_imm, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_info_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_inst_1_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_inst_1_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_jump_branch_info_jump_regiser, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_jump_branch_info_branch_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_executeStage_jump_branch_info_pred_branch, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_jump_branch_info_branch_target, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_executeStage_jump_branch_info_update_pht_index, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_valid, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_csr_in_pc, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [6:0]  io_csr_in_info_op, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_csr_in_info_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_csr_in_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_csr_out_rdata, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_csr_out_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_csr_out_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_csr_out_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input         io_csr_out_flush, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  input  [63:0] io_csr_out_target, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_bpu_pc, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [5:0]  io_bpu_update_pht_index, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_bpu_branch_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_bpu_branch, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_fetchUnit_flush, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_fetchUnit_target, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_decodeUnit_forward_0_exe_wen, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [4:0]  io_decodeUnit_forward_0_exe_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_decodeUnit_forward_0_exe_wdata, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_decodeUnit_forward_0_is_load, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_decodeUnit_forward_1_exe_wen, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [4:0]  io_decodeUnit_forward_1_exe_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_decodeUnit_forward_1_exe_wdata, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_decodeUnit_forward_1_is_load, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_pc, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_info_valid, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [2:0]  io_memoryStage_inst_0_info_fusel, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [6:0]  io_memoryStage_inst_0_info_op, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [4:0]  io_memoryStage_inst_0_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_info_imm, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_info_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_rd_info_wdata_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_rd_info_wdata_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_0_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_0_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_pc, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_info_valid, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [2:0]  io_memoryStage_inst_1_info_fusel, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [6:0]  io_memoryStage_inst_1_info_op, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_info_reg_wen, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [4:0]  io_memoryStage_inst_1_info_reg_waddr, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_info_imm, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_info_inst, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_rd_info_wdata_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_rd_info_wdata_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_src_info_src1_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_src_info_src2_data, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_exception_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_3, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_4, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_5, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_6, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_7, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_8, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_9, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_10, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output        io_memoryStage_inst_1_ex_interrupt_11, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_ex_tval_0, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_ex_tval_1, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_ex_tval_2, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_memoryStage_inst_1_ex_tval_12, // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
  output [63:0] io_dataMemory_addr // @[playground/src/pipeline/execute/ExecuteUnit.scala 13:14]
);
  wire  Fu_clock; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_reset; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_ctrl_allow_to_go; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_ctrl_stall; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_0_pc; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [2:0] Fu_io_inst_0_info_fusel; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [6:0] Fu_io_inst_0_info_op; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_0_info_imm; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_0_result_mdu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_0_result_alu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [2:0] Fu_io_inst_1_info_fusel; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [6:0] Fu_io_inst_1_info_op; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_1_info_imm; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_1_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_1_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_1_result_mdu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_inst_1_result_alu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_dataMemory_addr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_branch_pred_branch; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_branch_jump_regiser; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_branch_branch_target; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_branch_branch; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  Fu_io_branch_flush; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire [63:0] Fu_io_branch_target; // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
  wire  valid_0 = io_executeStage_inst_0_info_valid & io_ctrl_allow_to_go; // @[playground/src/pipeline/execute/ExecuteUnit.scala 39:53]
  wire  valid_1 = io_executeStage_inst_1_info_valid & io_ctrl_allow_to_go; // @[playground/src/pipeline/execute/ExecuteUnit.scala 39:53]
  wire [7:0] is_csr_lo = {4'h0,io_executeStage_inst_0_ex_exception_3,io_executeStage_inst_0_ex_exception_2,
    io_executeStage_inst_0_ex_exception_1,io_executeStage_inst_0_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _is_csr_T_2 = {2'h0,1'h0,io_executeStage_inst_0_ex_exception_12,io_executeStage_inst_0_ex_exception_11,1'h0
    ,io_executeStage_inst_0_ex_exception_9,io_executeStage_inst_0_ex_exception_8,is_csr_lo}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] is_csr_lo_1 = {io_executeStage_inst_0_ex_interrupt_5,io_executeStage_inst_0_ex_interrupt_4,
    io_executeStage_inst_0_ex_interrupt_3,io_executeStage_inst_0_ex_interrupt_2,io_executeStage_inst_0_ex_interrupt_1,
    io_executeStage_inst_0_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _is_csr_T_4 = {io_executeStage_inst_0_ex_interrupt_11,io_executeStage_inst_0_ex_interrupt_10,
    io_executeStage_inst_0_ex_interrupt_9,io_executeStage_inst_0_ex_interrupt_8,io_executeStage_inst_0_ex_interrupt_7,
    io_executeStage_inst_0_ex_interrupt_6,is_csr_lo_1}; // @[playground/src/defines/Util.scala 8:45]
  wire  _is_csr_T_6 = |_is_csr_T_2 | |_is_csr_T_4; // @[playground/src/defines/Util.scala 8:29]
  wire  is_csr_0 = io_executeStage_inst_0_info_fusel == 3'h3 & valid_0 & ~_is_csr_T_6; // @[playground/src/pipeline/execute/ExecuteUnit.scala 51:43]
  wire [7:0] is_csr_lo_2 = {4'h0,io_executeStage_inst_1_ex_exception_3,io_executeStage_inst_1_ex_exception_2,
    io_executeStage_inst_1_ex_exception_1,io_executeStage_inst_1_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _is_csr_T_11 = {2'h0,1'h0,io_executeStage_inst_1_ex_exception_12,io_executeStage_inst_1_ex_exception_11,1'h0
    ,io_executeStage_inst_1_ex_exception_9,io_executeStage_inst_1_ex_exception_8,is_csr_lo_2}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] is_csr_lo_3 = {io_executeStage_inst_1_ex_interrupt_5,io_executeStage_inst_1_ex_interrupt_4,
    io_executeStage_inst_1_ex_interrupt_3,io_executeStage_inst_1_ex_interrupt_2,io_executeStage_inst_1_ex_interrupt_1,
    io_executeStage_inst_1_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _is_csr_T_13 = {io_executeStage_inst_1_ex_interrupt_11,io_executeStage_inst_1_ex_interrupt_10,
    io_executeStage_inst_1_ex_interrupt_9,io_executeStage_inst_1_ex_interrupt_8,io_executeStage_inst_1_ex_interrupt_7,
    io_executeStage_inst_1_ex_interrupt_6,is_csr_lo_3}; // @[playground/src/defines/Util.scala 8:45]
  wire  _is_csr_T_15 = |_is_csr_T_11 | |_is_csr_T_13; // @[playground/src/defines/Util.scala 8:29]
  wire  is_csr_1 = io_executeStage_inst_1_info_fusel == 3'h3 & valid_1 & ~_is_csr_T_15; // @[playground/src/pipeline/execute/ExecuteUnit.scala 51:43]
  wire [1:0] _io_csr_in_valid_T = {is_csr_1,is_csr_0}; // @[playground/src/pipeline/execute/ExecuteUnit.scala 55:29]
  wire [63:0] _io_csr_in_pc_T = is_csr_0 ? io_executeStage_inst_0_pc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_pc_T_1 = is_csr_1 ? io_executeStage_inst_1_pc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_info_T = is_csr_0 ? io_executeStage_inst_0_info_inst : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_info_T_1 = is_csr_1 ? io_executeStage_inst_1_info_inst : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _io_csr_in_info_T_12 = is_csr_0 ? io_executeStage_inst_0_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _io_csr_in_info_T_13 = is_csr_1 ? io_executeStage_inst_1_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_src_info_T_3 = is_csr_0 ? io_executeStage_inst_0_src_info_src1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_src_info_T_4 = is_csr_1 ? io_executeStage_inst_1_src_info_src1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_3 = is_csr_0 ? io_executeStage_inst_0_ex_tval_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_4 = is_csr_1 ? io_executeStage_inst_1_ex_tval_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_36 = is_csr_0 ? io_executeStage_inst_0_ex_tval_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_37 = is_csr_1 ? io_executeStage_inst_1_ex_tval_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_memoryStage_inst_0_ex_T_5 = _is_csr_T_6 & io_executeStage_inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 98:47]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_1 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_1 : io_executeStage_inst_0_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_2 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_2 : io_executeStage_inst_0_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_3 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_3 : io_executeStage_inst_0_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_8 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_8 : io_executeStage_inst_0_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_9 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_9 : io_executeStage_inst_0_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_11 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_11 : io_executeStage_inst_0_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_exception_12 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_exception_12 : io_executeStage_inst_0_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_0 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_0 : io_executeStage_inst_0_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_1 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_1 : io_executeStage_inst_0_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_2 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_2 : io_executeStage_inst_0_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_3 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_3 : io_executeStage_inst_0_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_4 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_4 : io_executeStage_inst_0_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_5 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_5 : io_executeStage_inst_0_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_6 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_6 : io_executeStage_inst_0_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_7 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_7 : io_executeStage_inst_0_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_8 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_8 : io_executeStage_inst_0_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_9 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_9 : io_executeStage_inst_0_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_10 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_10 : io_executeStage_inst_0_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_T_7_interrupt_11 = 3'h3 == io_executeStage_inst_0_info_fusel ?
    io_csr_out_ex_interrupt_11 : io_executeStage_inst_0_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _io_memoryStage_inst_0_ex_T_7_tval_1 = 3'h3 == io_executeStage_inst_0_info_fusel ? io_csr_out_ex_tval_1 :
    io_executeStage_inst_0_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _io_memoryStage_inst_0_ex_T_7_tval_2 = 3'h3 == io_executeStage_inst_0_info_fusel ? io_csr_out_ex_tval_2 :
    io_executeStage_inst_0_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _io_memoryStage_inst_0_ex_T_7_tval_12 = 3'h3 == io_executeStage_inst_0_info_fusel ? io_csr_out_ex_tval_12
     : io_executeStage_inst_0_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_0_ex_exception_0_T_2 = io_fetchUnit_flush & |io_fetchUnit_target[1:0]; // @[playground/src/pipeline/execute/ExecuteUnit.scala 108:26]
  wire [63:0] _GEN_1 = 3'h1 == io_memoryStage_inst_0_info_fusel ? io_memoryStage_inst_0_rd_info_wdata_1 :
    io_memoryStage_inst_0_rd_info_wdata_0; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire [63:0] _GEN_2 = 3'h2 == io_memoryStage_inst_0_info_fusel ? io_memoryStage_inst_0_rd_info_wdata_2 : _GEN_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire [63:0] _GEN_3 = 3'h3 == io_memoryStage_inst_0_info_fusel ? io_memoryStage_inst_0_rd_info_wdata_3 : _GEN_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire [63:0] _GEN_4 = 3'h4 == io_memoryStage_inst_0_info_fusel ? io_memoryStage_inst_0_rd_info_wdata_4 : _GEN_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire  _io_memoryStage_inst_1_ex_T_5 = _is_csr_T_15 & io_executeStage_inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 98:47]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_1 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_1 : io_executeStage_inst_1_ex_exception_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_2 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_2 : io_executeStage_inst_1_ex_exception_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_3 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_3 : io_executeStage_inst_1_ex_exception_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_8 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_8 : io_executeStage_inst_1_ex_exception_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_9 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_9 : io_executeStage_inst_1_ex_exception_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_11 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_11 : io_executeStage_inst_1_ex_exception_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_exception_12 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_exception_12 : io_executeStage_inst_1_ex_exception_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_0 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_0 : io_executeStage_inst_1_ex_interrupt_0; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_1 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_1 : io_executeStage_inst_1_ex_interrupt_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_2 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_2 : io_executeStage_inst_1_ex_interrupt_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_3 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_3 : io_executeStage_inst_1_ex_interrupt_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_4 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_4 : io_executeStage_inst_1_ex_interrupt_4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_5 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_5 : io_executeStage_inst_1_ex_interrupt_5; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_6 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_6 : io_executeStage_inst_1_ex_interrupt_6; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_7 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_7 : io_executeStage_inst_1_ex_interrupt_7; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_8 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_8 : io_executeStage_inst_1_ex_interrupt_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_9 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_9 : io_executeStage_inst_1_ex_interrupt_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_10 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_10 : io_executeStage_inst_1_ex_interrupt_10; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire  _io_memoryStage_inst_1_ex_T_7_interrupt_11 = 3'h3 == io_executeStage_inst_1_info_fusel ?
    io_csr_out_ex_interrupt_11 : io_executeStage_inst_1_ex_interrupt_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _io_memoryStage_inst_1_ex_T_7_tval_1 = 3'h3 == io_executeStage_inst_1_info_fusel ? io_csr_out_ex_tval_1 :
    io_executeStage_inst_1_ex_tval_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _io_memoryStage_inst_1_ex_T_7_tval_2 = 3'h3 == io_executeStage_inst_1_info_fusel ? io_csr_out_ex_tval_2 :
    io_executeStage_inst_1_ex_tval_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _io_memoryStage_inst_1_ex_T_7_tval_12 = 3'h3 == io_executeStage_inst_1_info_fusel ? io_csr_out_ex_tval_12
     : io_executeStage_inst_1_ex_tval_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 100:80]
  wire [63:0] _GEN_7 = 3'h1 == io_memoryStage_inst_1_info_fusel ? io_memoryStage_inst_1_rd_info_wdata_1 :
    io_memoryStage_inst_1_rd_info_wdata_0; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire [63:0] _GEN_8 = 3'h2 == io_memoryStage_inst_1_info_fusel ? io_memoryStage_inst_1_rd_info_wdata_2 : _GEN_7; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire [63:0] _GEN_9 = 3'h3 == io_memoryStage_inst_1_info_fusel ? io_memoryStage_inst_1_rd_info_wdata_3 : _GEN_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  wire [63:0] _GEN_10 = 3'h4 == io_memoryStage_inst_1_info_fusel ? io_memoryStage_inst_1_rd_info_wdata_4 : _GEN_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  Fu Fu ( // @[playground/src/pipeline/execute/ExecuteUnit.scala 67:18]
    .clock(Fu_clock),
    .reset(Fu_reset),
    .io_ctrl_allow_to_go(Fu_io_ctrl_allow_to_go),
    .io_ctrl_stall(Fu_io_ctrl_stall),
    .io_inst_0_pc(Fu_io_inst_0_pc),
    .io_inst_0_info_valid(Fu_io_inst_0_info_valid),
    .io_inst_0_info_fusel(Fu_io_inst_0_info_fusel),
    .io_inst_0_info_op(Fu_io_inst_0_info_op),
    .io_inst_0_info_imm(Fu_io_inst_0_info_imm),
    .io_inst_0_src_info_src1_data(Fu_io_inst_0_src_info_src1_data),
    .io_inst_0_src_info_src2_data(Fu_io_inst_0_src_info_src2_data),
    .io_inst_0_result_mdu(Fu_io_inst_0_result_mdu),
    .io_inst_0_result_alu(Fu_io_inst_0_result_alu),
    .io_inst_1_info_valid(Fu_io_inst_1_info_valid),
    .io_inst_1_info_fusel(Fu_io_inst_1_info_fusel),
    .io_inst_1_info_op(Fu_io_inst_1_info_op),
    .io_inst_1_info_imm(Fu_io_inst_1_info_imm),
    .io_inst_1_src_info_src1_data(Fu_io_inst_1_src_info_src1_data),
    .io_inst_1_src_info_src2_data(Fu_io_inst_1_src_info_src2_data),
    .io_inst_1_result_mdu(Fu_io_inst_1_result_mdu),
    .io_inst_1_result_alu(Fu_io_inst_1_result_alu),
    .io_dataMemory_addr(Fu_io_dataMemory_addr),
    .io_branch_pred_branch(Fu_io_branch_pred_branch),
    .io_branch_jump_regiser(Fu_io_branch_jump_regiser),
    .io_branch_branch_target(Fu_io_branch_branch_target),
    .io_branch_branch(Fu_io_branch_branch),
    .io_branch_flush(Fu_io_branch_flush),
    .io_branch_target(Fu_io_branch_target)
  );
  assign io_ctrl_inst_0_is_load = io_executeStage_inst_0_info_fusel == 3'h1 & io_executeStage_inst_0_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteUnit.scala 45:57]
  assign io_ctrl_inst_0_reg_waddr = io_executeStage_inst_0_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 46:31]
  assign io_ctrl_inst_1_is_load = io_executeStage_inst_1_info_fusel == 3'h1 & io_executeStage_inst_1_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteUnit.scala 45:57]
  assign io_ctrl_inst_1_reg_waddr = io_executeStage_inst_1_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 46:31]
  assign io_ctrl_flush = io_fetchUnit_flush; // @[playground/src/pipeline/execute/ExecuteUnit.scala 42:17]
  assign io_ctrl_fu_stall = Fu_io_ctrl_stall; // @[playground/src/pipeline/execute/ExecuteUnit.scala 68:11]
  assign io_csr_in_valid = |_io_csr_in_valid_T; // @[playground/src/pipeline/execute/ExecuteUnit.scala 55:36]
  assign io_csr_in_pc = _io_csr_in_pc_T | _io_csr_in_pc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_info_op = _io_csr_in_info_T_12 | _io_csr_in_info_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_info_inst = _io_csr_in_info_T | _io_csr_in_info_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_src_info_src1_data = _io_csr_in_src_info_T_3 | _io_csr_in_src_info_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_1 = is_csr_0 & io_executeStage_inst_0_ex_exception_1 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_2 = is_csr_0 & io_executeStage_inst_0_ex_exception_2 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_3 = is_csr_0 & io_executeStage_inst_0_ex_exception_3 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_8 = is_csr_0 & io_executeStage_inst_0_ex_exception_8 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_9 = is_csr_0 & io_executeStage_inst_0_ex_exception_9 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_11 = is_csr_0 & io_executeStage_inst_0_ex_exception_11 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_exception_12 = is_csr_0 & io_executeStage_inst_0_ex_exception_12 | is_csr_1 &
    io_executeStage_inst_1_ex_exception_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_0 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_0 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_1 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_1 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_2 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_2 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_3 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_3 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_4 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_4 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_5 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_5 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_6 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_6 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_7 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_7 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_8 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_8 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_9 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_9 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_10 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_10 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_interrupt_11 = is_csr_0 & io_executeStage_inst_0_ex_interrupt_11 | is_csr_1 &
    io_executeStage_inst_1_ex_interrupt_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_tval_1 = _io_csr_in_ex_T_3 | _io_csr_in_ex_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_csr_in_ex_tval_12 = _io_csr_in_ex_T_36 | _io_csr_in_ex_T_37; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_bpu_pc = io_executeStage_inst_0_pc; // @[playground/src/pipeline/execute/ExecuteUnit.scala 80:27]
  assign io_bpu_update_pht_index = io_executeStage_jump_branch_info_update_pht_index[5:0]; // @[playground/src/pipeline/execute/ExecuteUnit.scala 81:27]
  assign io_bpu_branch_inst = io_executeStage_jump_branch_info_branch_inst; // @[playground/src/pipeline/execute/ExecuteUnit.scala 83:27]
  assign io_bpu_branch = Fu_io_branch_branch; // @[playground/src/pipeline/execute/ExecuteUnit.scala 82:27]
  assign io_fetchUnit_flush = valid_0 & io_ctrl_allow_to_go & (Fu_io_branch_flush | io_csr_out_flush); // @[playground/src/pipeline/execute/ExecuteUnit.scala 85:58]
  assign io_fetchUnit_target = io_csr_out_flush ? io_csr_out_target : Fu_io_branch_target; // @[playground/src/pipeline/execute/ExecuteUnit.scala 86:29]
  assign io_decodeUnit_forward_0_exe_wen = io_memoryStage_inst_0_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteUnit.scala 115:40]
  assign io_decodeUnit_forward_0_exe_waddr = io_memoryStage_inst_0_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 116:40]
  assign io_decodeUnit_forward_0_exe_wdata = 3'h5 == io_memoryStage_inst_0_info_fusel ?
    io_memoryStage_inst_0_rd_info_wdata_5 : _GEN_4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  assign io_decodeUnit_forward_0_is_load = io_ctrl_inst_0_is_load; // @[playground/src/pipeline/execute/ExecuteUnit.scala 118:40]
  assign io_decodeUnit_forward_1_exe_wen = io_memoryStage_inst_1_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteUnit.scala 115:40]
  assign io_decodeUnit_forward_1_exe_waddr = io_memoryStage_inst_1_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 116:40]
  assign io_decodeUnit_forward_1_exe_wdata = 3'h5 == io_memoryStage_inst_1_info_fusel ?
    io_memoryStage_inst_1_rd_info_wdata_5 : _GEN_10; // @[playground/src/pipeline/execute/ExecuteUnit.scala 117:{40,40}]
  assign io_decodeUnit_forward_1_is_load = io_ctrl_inst_1_is_load; // @[playground/src/pipeline/execute/ExecuteUnit.scala 118:40]
  assign io_memoryStage_inst_0_pc = io_executeStage_inst_0_pc; // @[playground/src/pipeline/execute/ExecuteUnit.scala 89:54]
  assign io_memoryStage_inst_0_info_valid = io_executeStage_inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_info_fusel = io_executeStage_inst_0_info_fusel; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_info_op = io_executeStage_inst_0_info_op; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_info_reg_wen = io_executeStage_inst_0_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_info_reg_waddr = io_executeStage_inst_0_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_info_imm = io_executeStage_inst_0_info_imm; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_info_inst = io_executeStage_inst_0_info_inst; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_0_rd_info_wdata_0 = Fu_io_inst_0_result_alu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 93:54]
  assign io_memoryStage_inst_0_rd_info_wdata_1 = 64'h0;
  assign io_memoryStage_inst_0_rd_info_wdata_2 = Fu_io_inst_0_result_mdu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 95:54]
  assign io_memoryStage_inst_0_rd_info_wdata_3 = io_csr_out_rdata; // @[playground/src/pipeline/execute/ExecuteUnit.scala 96:54]
  assign io_memoryStage_inst_0_rd_info_wdata_4 = 64'h0;
  assign io_memoryStage_inst_0_rd_info_wdata_5 = io_executeStage_inst_0_pc + 64'h4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 94:84]
  assign io_memoryStage_inst_0_src_info_src1_data = io_executeStage_inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 91:54]
  assign io_memoryStage_inst_0_src_info_src2_data = io_executeStage_inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 91:54]
  assign io_memoryStage_inst_0_ex_exception_0 = io_executeStage_inst_0_ex_exception_0 |
    _io_memoryStage_inst_0_ex_exception_0_T_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 107:64]
  assign io_memoryStage_inst_0_ex_exception_1 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_1 :
    _io_memoryStage_inst_0_ex_T_7_exception_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_exception_2 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_2 :
    _io_memoryStage_inst_0_ex_T_7_exception_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_exception_3 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_3 :
    _io_memoryStage_inst_0_ex_T_7_exception_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_exception_8 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_8 :
    _io_memoryStage_inst_0_ex_T_7_exception_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_exception_9 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_9 :
    _io_memoryStage_inst_0_ex_T_7_exception_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_exception_11 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_11
     : _io_memoryStage_inst_0_ex_T_7_exception_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_exception_12 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_exception_12
     : _io_memoryStage_inst_0_ex_T_7_exception_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_0 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_0 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_0; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_1 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_1 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_2 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_2 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_3 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_3 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_4 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_4 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_5 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_5 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_5; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_6 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_6 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_6; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_7 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_7 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_7; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_8 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_8 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_9 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_9 :
    _io_memoryStage_inst_0_ex_T_7_interrupt_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_10 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_10
     : _io_memoryStage_inst_0_ex_T_7_interrupt_10; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_interrupt_11 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_interrupt_11
     : _io_memoryStage_inst_0_ex_T_7_interrupt_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_tval_0 = io_executeStage_inst_0_ex_exception_0 ? io_executeStage_inst_0_ex_tval_0 :
    io_fetchUnit_target; // @[playground/src/pipeline/execute/ExecuteUnit.scala 109:62]
  assign io_memoryStage_inst_0_ex_tval_1 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_tval_1 :
    _io_memoryStage_inst_0_ex_T_7_tval_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_tval_2 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_tval_2 :
    _io_memoryStage_inst_0_ex_T_7_tval_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_0_ex_tval_12 = _io_memoryStage_inst_0_ex_T_5 ? io_executeStage_inst_0_ex_tval_12 :
    _io_memoryStage_inst_0_ex_T_7_tval_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_pc = io_executeStage_inst_1_pc; // @[playground/src/pipeline/execute/ExecuteUnit.scala 89:54]
  assign io_memoryStage_inst_1_info_valid = io_executeStage_inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_info_fusel = io_executeStage_inst_1_info_fusel; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_info_op = io_executeStage_inst_1_info_op; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_info_reg_wen = io_executeStage_inst_1_info_reg_wen; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_info_reg_waddr = io_executeStage_inst_1_info_reg_waddr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_info_imm = io_executeStage_inst_1_info_imm; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_info_inst = io_executeStage_inst_1_info_inst; // @[playground/src/pipeline/execute/ExecuteUnit.scala 90:54]
  assign io_memoryStage_inst_1_rd_info_wdata_0 = Fu_io_inst_1_result_alu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 93:54]
  assign io_memoryStage_inst_1_rd_info_wdata_1 = 64'h0;
  assign io_memoryStage_inst_1_rd_info_wdata_2 = Fu_io_inst_1_result_mdu; // @[playground/src/pipeline/execute/ExecuteUnit.scala 95:54]
  assign io_memoryStage_inst_1_rd_info_wdata_3 = io_csr_out_rdata; // @[playground/src/pipeline/execute/ExecuteUnit.scala 96:54]
  assign io_memoryStage_inst_1_rd_info_wdata_4 = 64'h0;
  assign io_memoryStage_inst_1_rd_info_wdata_5 = io_executeStage_inst_1_pc + 64'h4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 94:84]
  assign io_memoryStage_inst_1_src_info_src1_data = io_executeStage_inst_1_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 91:54]
  assign io_memoryStage_inst_1_src_info_src2_data = io_executeStage_inst_1_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 91:54]
  assign io_memoryStage_inst_1_ex_exception_0 = io_executeStage_inst_1_ex_exception_0 |
    _io_memoryStage_inst_0_ex_exception_0_T_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 107:64]
  assign io_memoryStage_inst_1_ex_exception_1 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_1 :
    _io_memoryStage_inst_1_ex_T_7_exception_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_exception_2 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_2 :
    _io_memoryStage_inst_1_ex_T_7_exception_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_exception_3 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_3 :
    _io_memoryStage_inst_1_ex_T_7_exception_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_exception_8 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_8 :
    _io_memoryStage_inst_1_ex_T_7_exception_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_exception_9 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_9 :
    _io_memoryStage_inst_1_ex_T_7_exception_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_exception_11 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_11
     : _io_memoryStage_inst_1_ex_T_7_exception_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_exception_12 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_exception_12
     : _io_memoryStage_inst_1_ex_T_7_exception_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_0 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_0 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_0; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_1 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_1 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_2 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_2 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_3 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_3 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_3; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_4 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_4 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_4; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_5 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_5 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_5; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_6 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_6 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_6; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_7 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_7 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_7; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_8 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_8 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_8; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_9 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_9 :
    _io_memoryStage_inst_1_ex_T_7_interrupt_9; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_10 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_10
     : _io_memoryStage_inst_1_ex_T_7_interrupt_10; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_interrupt_11 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_interrupt_11
     : _io_memoryStage_inst_1_ex_T_7_interrupt_11; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_tval_0 = io_executeStage_inst_1_ex_exception_0 ? io_executeStage_inst_1_ex_tval_0 :
    io_fetchUnit_target; // @[playground/src/pipeline/execute/ExecuteUnit.scala 109:62]
  assign io_memoryStage_inst_1_ex_tval_1 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_tval_1 :
    _io_memoryStage_inst_1_ex_T_7_tval_1; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_tval_2 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_tval_2 :
    _io_memoryStage_inst_1_ex_T_7_tval_2; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_memoryStage_inst_1_ex_tval_12 = _io_memoryStage_inst_1_ex_T_5 ? io_executeStage_inst_1_ex_tval_12 :
    _io_memoryStage_inst_1_ex_T_7_tval_12; // @[playground/src/pipeline/execute/ExecuteUnit.scala 97:37]
  assign io_dataMemory_addr = Fu_io_dataMemory_addr; // @[playground/src/pipeline/execute/ExecuteUnit.scala 78:22]
  assign Fu_clock = clock;
  assign Fu_reset = reset;
  assign Fu_io_ctrl_allow_to_go = io_ctrl_fu_allow_to_go; // @[playground/src/pipeline/execute/ExecuteUnit.scala 68:11]
  assign Fu_io_inst_0_pc = io_executeStage_inst_0_pc; // @[playground/src/pipeline/execute/ExecuteUnit.scala 70:25]
  assign Fu_io_inst_0_info_valid = io_executeStage_inst_0_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_0_info_fusel = io_executeStage_inst_0_info_fusel; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_0_info_op = io_executeStage_inst_0_info_op; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_0_info_imm = io_executeStage_inst_0_info_imm; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_0_src_info_src1_data = io_executeStage_inst_0_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 72:25]
  assign Fu_io_inst_0_src_info_src2_data = io_executeStage_inst_0_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 72:25]
  assign Fu_io_inst_1_info_valid = io_executeStage_inst_1_info_valid; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_1_info_fusel = io_executeStage_inst_1_info_fusel; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_1_info_op = io_executeStage_inst_1_info_op; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_1_info_imm = io_executeStage_inst_1_info_imm; // @[playground/src/pipeline/execute/ExecuteUnit.scala 71:25]
  assign Fu_io_inst_1_src_info_src1_data = io_executeStage_inst_1_src_info_src1_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 72:25]
  assign Fu_io_inst_1_src_info_src2_data = io_executeStage_inst_1_src_info_src2_data; // @[playground/src/pipeline/execute/ExecuteUnit.scala 72:25]
  assign Fu_io_branch_pred_branch = io_executeStage_jump_branch_info_pred_branch; // @[playground/src/pipeline/execute/ExecuteUnit.scala 74:27]
  assign Fu_io_branch_jump_regiser = io_executeStage_jump_branch_info_jump_regiser; // @[playground/src/pipeline/execute/ExecuteUnit.scala 75:27]
  assign Fu_io_branch_branch_target = io_executeStage_jump_branch_info_branch_target; // @[playground/src/pipeline/execute/ExecuteUnit.scala 76:27]
endmodule
module Csr(
  input         clock,
  input         reset,
  input         io_ext_int_ei, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_ext_int_ti, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_ext_int_si, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [1:0]  io_decodeUnit_mode, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [11:0] io_decodeUnit_interrupt, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_valid, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_executeUnit_in_pc, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [6:0]  io_executeUnit_in_info_op, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_executeUnit_in_info_inst, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_executeUnit_in_src_info_src1_data, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_exception_12, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_0, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_4, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_5, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_6, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_7, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_10, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_executeUnit_in_ex_interrupt_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_executeUnit_in_ex_tval_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_executeUnit_in_ex_tval_12, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_executeUnit_out_rdata, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_exception_12, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_0, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_4, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_5, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_6, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_7, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_10, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_ex_interrupt_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_executeUnit_out_ex_tval_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_executeUnit_out_ex_tval_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_executeUnit_out_ex_tval_12, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_executeUnit_out_flush, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_executeUnit_out_target, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_pc, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_0, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_4, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_5, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_6, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_7, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_10, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_12, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_13, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_14, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_exception_15, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_0, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_4, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_5, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_6, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_7, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_10, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_ex_interrupt_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_0, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_1, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_2, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_3, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_4, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_5, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_6, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_7, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_8, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_9, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_10, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_11, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_12, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_13, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_14, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_ex_tval_15, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_info_valid, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [2:0]  io_memoryUnit_in_info_fusel, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [6:0]  io_memoryUnit_in_info_op, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_lr_wen, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input         io_memoryUnit_in_lr_wbit, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  input  [63:0] io_memoryUnit_in_lr_waddr, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_memoryUnit_out_flush, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_memoryUnit_out_target, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output        io_memoryUnit_out_lr, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_memoryUnit_out_lr_addr, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_tlb_satp, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [63:0] io_tlb_mstatus, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [1:0]  io_tlb_imode, // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
  output [1:0]  io_tlb_dmode // @[playground/src/pipeline/execute/fu/Csr.scala 58:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mstatus; // @[playground/src/pipeline/execute/fu/Csr.scala 81:26]
  reg [63:0] medeleg; // @[playground/src/pipeline/execute/fu/Csr.scala 93:27]
  reg [63:0] mideleg; // @[playground/src/pipeline/execute/fu/Csr.scala 94:27]
  reg [63:0] mie; // @[playground/src/pipeline/execute/fu/Csr.scala 95:27]
  reg [63:0] mtvec; // @[playground/src/pipeline/execute/fu/Csr.scala 96:27]
  reg [63:0] mcounteren; // @[playground/src/pipeline/execute/fu/Csr.scala 97:27]
  reg [63:0] mscratch; // @[playground/src/pipeline/execute/fu/Csr.scala 100:27]
  reg [63:0] mepc; // @[playground/src/pipeline/execute/fu/Csr.scala 101:27]
  reg [63:0] mcause; // @[playground/src/pipeline/execute/fu/Csr.scala 102:27]
  reg [63:0] mtval; // @[playground/src/pipeline/execute/fu/Csr.scala 103:27]
  reg [63:0] mipReg; // @[playground/src/pipeline/execute/fu/Csr.scala 105:27]
  wire [11:0] _mip_T = {io_ext_int_ei,1'h0,1'h0,1'h0,io_ext_int_ti,1'h0,2'h0,io_ext_int_si,3'h0}; // @[playground/src/pipeline/execute/fu/Csr.scala 107:28]
  wire [63:0] _GEN_77 = {{52'd0}, _mip_T}; // @[playground/src/pipeline/execute/fu/Csr.scala 107:35]
  wire [63:0] mip = _GEN_77 | mipReg; // @[playground/src/pipeline/execute/fu/Csr.scala 107:35]
  reg [63:0] mcycle; // @[playground/src/pipeline/execute/fu/Csr.scala 122:23]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[playground/src/pipeline/execute/fu/Csr.scala 123:20]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[playground/src/pipeline/execute/fu/Csr.scala 133:35]
  reg [63:0] stvec; // @[playground/src/pipeline/execute/fu/Csr.scala 134:27]
  reg [63:0] scounteren; // @[playground/src/pipeline/execute/fu/Csr.scala 135:27]
  reg [63:0] sscratch; // @[playground/src/pipeline/execute/fu/Csr.scala 138:25]
  reg [63:0] sepc; // @[playground/src/pipeline/execute/fu/Csr.scala 139:25]
  reg [63:0] scause; // @[playground/src/pipeline/execute/fu/Csr.scala 140:25]
  reg [63:0] stval; // @[playground/src/pipeline/execute/fu/Csr.scala 141:25]
  reg [63:0] satp; // @[playground/src/pipeline/execute/fu/Csr.scala 146:21]
  reg  lr; // @[playground/src/pipeline/execute/fu/Csr.scala 159:25]
  reg [63:0] lr_addr; // @[playground/src/pipeline/execute/fu/Csr.scala 160:25]
  wire  _wdata_T_6 = 7'h1 == io_executeUnit_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _wdata_T_12 = _wdata_T_6 ? io_executeUnit_in_src_info_src1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wdata_T_7 = 7'h2 == io_executeUnit_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [11:0] addr = io_executeUnit_in_info_inst[31:20]; // @[playground/src/pipeline/execute/fu/Csr.scala 276:42]
  wire  _rdata_T_29 = 12'h180 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_58 = _rdata_T_29 ? satp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_30 = 12'h140 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_59 = _rdata_T_30 ? sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_87 = _rdata_T_58 | _rdata_T_59; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_31 = 12'h306 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_60 = _rdata_T_31 ? mcounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_88 = _rdata_T_87 | _rdata_T_60; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_32 = 12'hf11 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_T_33 = 12'h104 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_4 = mie & sieMask; // @[playground/src/defines/Util.scala 112:84]
  wire [63:0] _rdata_T_62 = _rdata_T_33 ? _rdata_T_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_90 = _rdata_T_88 | _rdata_T_62; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_34 = 12'h144 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_5 = mip & sieMask; // @[playground/src/defines/Util.scala 112:84]
  wire [63:0] _rdata_T_63 = _rdata_T_34 ? _rdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_91 = _rdata_T_90 | _rdata_T_63; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_35 = 12'h7a1 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_T_36 = 12'h100 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_7 = mstatus & 64'h80000003000de762; // @[playground/src/defines/Util.scala 112:84]
  wire [63:0] _rdata_T_65 = _rdata_T_36 ? _rdata_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_93 = _rdata_T_91 | _rdata_T_65; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_37 = 12'h305 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_66 = _rdata_T_37 ? mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_94 = _rdata_T_93 | _rdata_T_66; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_38 = 12'h304 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_67 = _rdata_T_38 ? mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_95 = _rdata_T_94 | _rdata_T_67; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_39 = 12'h300 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_68 = _rdata_T_39 ? mstatus : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_96 = _rdata_T_95 | _rdata_T_68; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_40 = 12'h344 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_69 = _rdata_T_40 ? mip : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_97 = _rdata_T_96 | _rdata_T_69; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_41 = 12'h303 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_70 = _rdata_T_41 ? mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_98 = _rdata_T_97 | _rdata_T_70; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_42 = 12'hf13 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_T_43 = 12'h340 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_72 = _rdata_T_43 ? mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_100 = _rdata_T_98 | _rdata_T_72; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_44 = 12'h142 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_73 = _rdata_T_44 ? scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_101 = _rdata_T_100 | _rdata_T_73; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_45 = 12'hc00 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_74 = _rdata_T_45 ? mcycle : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_102 = _rdata_T_101 | _rdata_T_74; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_46 = 12'hf12 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_T_47 = 12'h302 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_76 = _rdata_T_47 ? medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_104 = _rdata_T_102 | _rdata_T_76; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_48 = 12'h105 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_77 = _rdata_T_48 ? stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_105 = _rdata_T_104 | _rdata_T_77; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_49 = 12'h141 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_78 = _rdata_T_49 ? sepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_106 = _rdata_T_105 | _rdata_T_78; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_50 = 12'h342 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_79 = _rdata_T_50 ? mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_107 = _rdata_T_106 | _rdata_T_79; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_51 = 12'h143 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_80 = _rdata_T_51 ? stval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_108 = _rdata_T_107 | _rdata_T_80; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_52 = 12'h301 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_81 = _rdata_T_52 ? 64'h8000000000141101 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_109 = _rdata_T_108 | _rdata_T_81; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_53 = 12'h7a0 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_82 = _rdata_T_53 ? 64'h1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_110 = _rdata_T_109 | _rdata_T_82; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_54 = 12'hf14 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_T_55 = 12'h341 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_84 = _rdata_T_55 ? mepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_112 = _rdata_T_110 | _rdata_T_84; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_56 = 12'h343 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_85 = _rdata_T_56 ? mtval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_113 = _rdata_T_112 | _rdata_T_85; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_57 = 12'h106 == addr; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_T_86 = _rdata_T_57 ? scounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T = rdata | io_executeUnit_in_src_info_src1_data; // @[playground/src/pipeline/execute/fu/Csr.scala 283:34]
  wire [63:0] _wdata_T_13 = _wdata_T_7 ? _wdata_T : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_18 = _wdata_T_12 | _wdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wdata_T_8 = 7'h3 == io_executeUnit_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _wdata_T_1 = ~io_executeUnit_in_src_info_src1_data; // @[playground/src/pipeline/execute/fu/Csr.scala 284:36]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[playground/src/pipeline/execute/fu/Csr.scala 284:34]
  wire [63:0] _wdata_T_14 = _wdata_T_8 ? _wdata_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_19 = _wdata_T_18 | _wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wdata_T_9 = 7'h5 == io_executeUnit_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] csri = {59'h0,io_executeUnit_in_info_inst[19:15]}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _wdata_T_15 = _wdata_T_9 ? csri : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_20 = _wdata_T_19 | _wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wdata_T_10 = 7'h6 == io_executeUnit_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _wdata_T_3 = rdata | csri; // @[playground/src/pipeline/execute/fu/Csr.scala 286:34]
  wire [63:0] _wdata_T_16 = _wdata_T_10 ? _wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_21 = _wdata_T_20 | _wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wdata_T_11 = 7'h7 == io_executeUnit_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _wdata_T_4 = ~csri; // @[playground/src/pipeline/execute/fu/Csr.scala 287:36]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[playground/src/pipeline/execute/fu/Csr.scala 287:34]
  wire [63:0] _wdata_T_17 = _wdata_T_11 ? _wdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] wdata = _wdata_T_21 | _wdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _mstatus_wmask_T_29 = 2'h3 == wdata[12:11] | 2'h1 == wdata[12:11] | 2'h0 == wdata[12:11]; // @[playground/src/pipeline/execute/fu/Csr.scala 178:42]
  wire [63:0] mstatus_wmask = _mstatus_wmask_T_29 ? 64'h7e19aa : 64'h7e01aa; // @[playground/src/pipeline/execute/fu/Csr.scala 177:26]
  reg [1:0] mode; // @[playground/src/pipeline/execute/fu/Csr.scala 234:21]
  wire  mip_raise_interrupt_s_u = mip[0]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_s_s = mip[1]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_s_h = mip[2]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_s_m = mip[3]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_t_u = mip[4]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_t_s = mip[5]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_t_h = mip[6]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_t_m = mip[7]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_e_u = mip[8]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_e_h = mip[10]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_e_m = mip[11]; // @[playground/src/pipeline/execute/fu/Csr.scala 244:50]
  wire  mip_raise_interrupt_e_s = mip[9] | io_ext_int_ei; // @[playground/src/pipeline/execute/fu/Csr.scala 245:62]
  wire  mstatusBundle_ie_u = mstatus[0]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_ie_s = mstatus[1]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_ie_h = mstatus[2]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_ie_m = mstatus[3]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_pie_u = mstatus[4]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_pie_s = mstatus[5]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_pie_h = mstatus[6]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_pie_m = mstatus[7]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_spp = mstatus[8]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [1:0] mstatusBundle_hpp = mstatus[10:9]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [1:0] mstatusBundle_mpp = mstatus[12:11]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [1:0] mstatusBundle_fs = mstatus[14:13]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [1:0] mstatusBundle_xs = mstatus[16:15]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_mprv = mstatus[17]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_sum = mstatus[18]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_mxr = mstatus[19]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_tvm = mstatus[20]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_tw = mstatus[21]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_tsr = mstatus[22]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [8:0] mstatusBundle_pad0 = mstatus[31:23]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [1:0] mstatusBundle_uxl = mstatus[33:32]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [1:0] mstatusBundle_sxl = mstatus[35:34]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [26:0] mstatusBundle_pad1 = mstatus[62:36]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire  mstatusBundle_sd = mstatus[63]; // @[playground/src/pipeline/execute/fu/Csr.scala 247:39]
  wire [5:0] ideleg_lo = {mip_raise_interrupt_t_s,mip_raise_interrupt_t_u,mip_raise_interrupt_s_m,
    mip_raise_interrupt_s_h,mip_raise_interrupt_s_s,mip_raise_interrupt_s_u}; // @[playground/src/pipeline/execute/fu/Csr.scala 249:47]
  wire [11:0] _ideleg_T = {mip_raise_interrupt_e_m,mip_raise_interrupt_e_h,mip_raise_interrupt_e_s,
    mip_raise_interrupt_e_u,mip_raise_interrupt_t_m,mip_raise_interrupt_t_h,ideleg_lo}; // @[playground/src/pipeline/execute/fu/Csr.scala 249:47]
  wire [63:0] _GEN_78 = {{52'd0}, _ideleg_T}; // @[playground/src/pipeline/execute/fu/Csr.scala 249:25]
  wire [63:0] ideleg = mideleg & _GEN_78; // @[playground/src/pipeline/execute/fu/Csr.scala 249:25]
  wire  _interrupt_enable_0_T_3 = mode == 2'h1 & mstatusBundle_ie_s | mode < 2'h1; // @[playground/src/pipeline/execute/fu/Csr.scala 252:46]
  wire  _interrupt_enable_0_T_6 = mode < 2'h3; // @[playground/src/pipeline/execute/fu/Csr.scala 253:55]
  wire  _interrupt_enable_0_T_7 = mode == 2'h3 & mstatusBundle_ie_m | mode < 2'h3; // @[playground/src/pipeline/execute/fu/Csr.scala 253:46]
  wire  interrupt_enable_0 = ideleg[0] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_1 = ideleg[1] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_2 = ideleg[2] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_3 = ideleg[3] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_4 = ideleg[4] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_5 = ideleg[5] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_6 = ideleg[6] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_7 = ideleg[7] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_8 = ideleg[8] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_9 = ideleg[9] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_10 = ideleg[10] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire  interrupt_enable_11 = ideleg[11] ? _interrupt_enable_0_T_3 : _interrupt_enable_0_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 250:51]
  wire [11:0] _io_decodeUnit_interrupt_T_2 = mie[11:0] & _ideleg_T; // @[playground/src/pipeline/execute/fu/Csr.scala 258:50]
  wire [5:0] io_decodeUnit_interrupt_lo_1 = {interrupt_enable_5,interrupt_enable_4,interrupt_enable_3,interrupt_enable_2
    ,interrupt_enable_1,interrupt_enable_0}; // @[playground/src/pipeline/execute/fu/Csr.scala 258:98]
  wire [11:0] _io_decodeUnit_interrupt_T_3 = {interrupt_enable_11,interrupt_enable_10,interrupt_enable_9,
    interrupt_enable_8,interrupt_enable_7,interrupt_enable_6,io_decodeUnit_interrupt_lo_1}; // @[playground/src/pipeline/execute/fu/Csr.scala 258:98]
  wire [7:0] raise_exception_lo = {io_memoryUnit_in_ex_exception_7,io_memoryUnit_in_ex_exception_6,
    io_memoryUnit_in_ex_exception_5,io_memoryUnit_in_ex_exception_4,io_memoryUnit_in_ex_exception_3,
    io_memoryUnit_in_ex_exception_2,io_memoryUnit_in_ex_exception_1,io_memoryUnit_in_ex_exception_0}; // @[playground/src/pipeline/execute/fu/Csr.scala 268:42]
  wire [15:0] _raise_exception_T = {io_memoryUnit_in_ex_exception_15,io_memoryUnit_in_ex_exception_14,
    io_memoryUnit_in_ex_exception_13,io_memoryUnit_in_ex_exception_12,io_memoryUnit_in_ex_exception_11,
    io_memoryUnit_in_ex_exception_10,io_memoryUnit_in_ex_exception_9,io_memoryUnit_in_ex_exception_8,raise_exception_lo}
    ; // @[playground/src/pipeline/execute/fu/Csr.scala 268:42]
  wire  raise_exception = |_raise_exception_T & io_memoryUnit_in_info_valid; // @[playground/src/pipeline/execute/fu/Csr.scala 268:53]
  wire [5:0] raise_interrupt_lo = {io_memoryUnit_in_ex_interrupt_5,io_memoryUnit_in_ex_interrupt_4,
    io_memoryUnit_in_ex_interrupt_3,io_memoryUnit_in_ex_interrupt_2,io_memoryUnit_in_ex_interrupt_1,
    io_memoryUnit_in_ex_interrupt_0}; // @[playground/src/pipeline/execute/fu/Csr.scala 269:42]
  wire [11:0] _raise_interrupt_T = {io_memoryUnit_in_ex_interrupt_11,io_memoryUnit_in_ex_interrupt_10,
    io_memoryUnit_in_ex_interrupt_9,io_memoryUnit_in_ex_interrupt_8,io_memoryUnit_in_ex_interrupt_7,
    io_memoryUnit_in_ex_interrupt_6,raise_interrupt_lo}; // @[playground/src/pipeline/execute/fu/Csr.scala 269:42]
  wire  raise_interrupt = |_raise_interrupt_T & io_memoryUnit_in_info_valid; // @[playground/src/pipeline/execute/fu/Csr.scala 269:53]
  wire  raise_exc_int = raise_exception | raise_interrupt; // @[playground/src/pipeline/execute/fu/Csr.scala 270:41]
  wire  valid = io_executeUnit_in_valid & ~io_memoryUnit_out_flush; // @[playground/src/pipeline/execute/fu/Csr.scala 272:39]
  wire  satp_legal = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[playground/src/pipeline/execute/fu/Csr.scala 291:62]
  wire  _write_T_1 = ~io_executeUnit_in_info_op[3]; // @[playground/src/defines/isa/Instructions.scala 159:27]
  wire  write = valid & _write_T_1 & (addr != 12'h180 | satp_legal); // @[playground/src/pipeline/execute/fu/Csr.scala 292:53]
  wire  only_read = (_wdata_T_7 | _wdata_T_10 | _wdata_T_8 | _wdata_T_11) & io_executeUnit_in_src_info_src1_data == 64'h0
    ; // @[playground/src/pipeline/execute/fu/Csr.scala 294:96]
  wire  illegal_mode = mode < addr[9:8]; // @[playground/src/pipeline/execute/fu/Csr.scala 295:29]
  wire  illegal_write = write & addr[11:10] == 2'h3 & ~only_read; // @[playground/src/pipeline/execute/fu/Csr.scala 296:60]
  wire  illegal_access = illegal_mode | illegal_write; // @[playground/src/pipeline/execute/fu/Csr.scala 297:37]
  wire  wen = write & ~illegal_access; // @[playground/src/pipeline/execute/fu/Csr.scala 298:30]
  wire  _T_105 = addr == 12'h180; // @[playground/src/defines/Util.scala 115:66]
  wire [63:0] _mie_T = wdata & sieMask; // @[playground/src/defines/Util.scala 58:14]
  wire [63:0] _mie_T_1 = ~sieMask; // @[playground/src/defines/Util.scala 58:39]
  wire [63:0] _mie_T_2 = mie & _mie_T_1; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _mie_T_3 = _mie_T | _mie_T_2; // @[playground/src/defines/Util.scala 58:26]
  wire [63:0] _mstatus_T_1 = wdata & 64'hc0122; // @[playground/src/defines/Util.scala 58:14]
  wire [63:0] _mstatus_T_3 = mstatus & 64'hfffffffffff3fedd; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _mstatus_T_4 = _mstatus_T_1 | _mstatus_T_3; // @[playground/src/defines/Util.scala 58:26]
  wire [1:0] mstatus_mstatusOld_fs = _mstatus_T_4[14:13]; // @[playground/src/pipeline/execute/fu/Csr.scala 172:47]
  wire [63:0] mstatus_mstatusNew = {mstatus_mstatusOld_fs == 2'h3,_mstatus_T_4[62:0]}; // @[playground/src/pipeline/execute/fu/Csr.scala 173:25]
  wire [63:0] _GEN_6 = wen & addr == 12'h100 ? mstatus_mstatusNew : mstatus; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 81:26]
  wire [63:0] _mstatus_T_5 = wdata & mstatus_wmask; // @[playground/src/defines/Util.scala 58:14]
  wire [63:0] _mstatus_T_6 = ~mstatus_wmask; // @[playground/src/defines/Util.scala 58:39]
  wire [63:0] _mstatus_T_7 = mstatus & _mstatus_T_6; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _mstatus_T_8 = _mstatus_T_5 | _mstatus_T_7; // @[playground/src/defines/Util.scala 58:26]
  wire [63:0] _GEN_9 = wen & addr == 12'h300 ? _mstatus_T_8 : _GEN_6; // @[playground/src/defines/Util.scala 115:{73,77}]
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[playground/src/defines/Util.scala 58:14]
  wire [63:0] _mideleg_T_2 = mideleg & 64'hfffffffffffffddd; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _mideleg_T_3 = _mideleg_T | _mideleg_T_2; // @[playground/src/defines/Util.scala 58:26]
  wire [63:0] _GEN_12 = wen & addr == 12'h142 ? wdata : scause; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 140:25]
  wire [63:0] _medeleg_T = wdata & 64'hbbff; // @[playground/src/defines/Util.scala 58:14]
  wire [63:0] _medeleg_T_2 = medeleg & 64'hffffffffffff4400; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[playground/src/defines/Util.scala 58:26]
  wire [63:0] _GEN_16 = wen & addr == 12'h141 ? wdata : sepc; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 139:25]
  wire [63:0] _GEN_17 = wen & addr == 12'h342 ? wdata : mcause; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 102:27]
  wire [63:0] _GEN_18 = wen & addr == 12'h143 ? wdata : stval; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 141:25]
  wire [63:0] _GEN_19 = wen & addr == 12'h341 ? wdata : mepc; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 101:27]
  wire [63:0] _GEN_20 = wen & addr == 12'h343 ? wdata : mtval; // @[playground/src/defines/Util.scala 115:{73,77} playground/src/pipeline/execute/fu/Csr.scala 103:27]
  wire  _illegal_addr_illegalAddr_T_1 = _rdata_T_29 ? 1'h0 : 1'h1; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_3 = _rdata_T_30 ? 1'h0 : _illegal_addr_illegalAddr_T_1; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_5 = _rdata_T_31 ? 1'h0 : _illegal_addr_illegalAddr_T_3; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_7 = _rdata_T_32 ? 1'h0 : _illegal_addr_illegalAddr_T_5; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_9 = _rdata_T_33 ? 1'h0 : _illegal_addr_illegalAddr_T_7; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_11 = _rdata_T_34 ? 1'h0 : _illegal_addr_illegalAddr_T_9; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_13 = _rdata_T_35 ? 1'h0 : _illegal_addr_illegalAddr_T_11; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_15 = _rdata_T_36 ? 1'h0 : _illegal_addr_illegalAddr_T_13; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_17 = _rdata_T_37 ? 1'h0 : _illegal_addr_illegalAddr_T_15; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_19 = _rdata_T_38 ? 1'h0 : _illegal_addr_illegalAddr_T_17; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_21 = _rdata_T_39 ? 1'h0 : _illegal_addr_illegalAddr_T_19; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_23 = _rdata_T_40 ? 1'h0 : _illegal_addr_illegalAddr_T_21; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_25 = _rdata_T_41 ? 1'h0 : _illegal_addr_illegalAddr_T_23; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_27 = _rdata_T_42 ? 1'h0 : _illegal_addr_illegalAddr_T_25; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_29 = _rdata_T_43 ? 1'h0 : _illegal_addr_illegalAddr_T_27; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_31 = _rdata_T_44 ? 1'h0 : _illegal_addr_illegalAddr_T_29; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_33 = _rdata_T_45 ? 1'h0 : _illegal_addr_illegalAddr_T_31; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_35 = _rdata_T_46 ? 1'h0 : _illegal_addr_illegalAddr_T_33; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_37 = _rdata_T_47 ? 1'h0 : _illegal_addr_illegalAddr_T_35; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_39 = _rdata_T_48 ? 1'h0 : _illegal_addr_illegalAddr_T_37; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_41 = _rdata_T_49 ? 1'h0 : _illegal_addr_illegalAddr_T_39; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_43 = _rdata_T_50 ? 1'h0 : _illegal_addr_illegalAddr_T_41; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_45 = _rdata_T_51 ? 1'h0 : _illegal_addr_illegalAddr_T_43; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_47 = _rdata_T_52 ? 1'h0 : _illegal_addr_illegalAddr_T_45; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_49 = _rdata_T_53 ? 1'h0 : _illegal_addr_illegalAddr_T_47; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_51 = _rdata_T_54 ? 1'h0 : _illegal_addr_illegalAddr_T_49; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_53 = _rdata_T_55 ? 1'h0 : _illegal_addr_illegalAddr_T_51; // @[playground/src/defines/Util.scala 51:28]
  wire  _illegal_addr_illegalAddr_T_55 = _rdata_T_56 ? 1'h0 : _illegal_addr_illegalAddr_T_53; // @[playground/src/defines/Util.scala 51:28]
  wire  illegal_addr = _rdata_T_57 ? 1'h0 : _illegal_addr_illegalAddr_T_55; // @[playground/src/defines/Util.scala 51:28]
  wire [63:0] _mipReg_T = wdata & 64'haaa; // @[playground/src/defines/Util.scala 58:14]
  wire [63:0] _mipReg_T_2 = mipReg & 64'hfffffffffffff555; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _mipReg_T_3 = _mipReg_T | _mipReg_T_2; // @[playground/src/defines/Util.scala 58:26]
  wire [63:0] _mipReg_T_6 = mipReg & _mie_T_1; // @[playground/src/defines/Util.scala 58:37]
  wire [63:0] _mipReg_T_7 = _mie_T | _mipReg_T_6; // @[playground/src/defines/Util.scala 58:26]
  wire  _isMret_T = io_memoryUnit_in_info_fusel == 3'h3; // @[playground/src/defines/Util.scala 14:16]
  wire  _isMret_T_2 = io_memoryUnit_in_info_fusel == 3'h3 & io_memoryUnit_in_info_op == 7'ha; // @[playground/src/defines/Util.scala 14:31]
  wire  isMret = _isMret_T_2 & io_memoryUnit_in_info_valid; // @[playground/src/pipeline/execute/fu/Csr.scala 312:38]
  wire  _isSret_T_2 = _isMret_T & io_memoryUnit_in_info_op == 7'hb; // @[playground/src/defines/Util.scala 20:31]
  wire  isSret = _isSret_T_2 & io_memoryUnit_in_info_valid; // @[playground/src/pipeline/execute/fu/Csr.scala 313:38]
  wire  ret = isMret | isSret; // @[playground/src/pipeline/execute/fu/Csr.scala 314:17]
  wire [2:0] _exceptionNO_T = io_memoryUnit_in_ex_exception_5 ? 3'h5 : 3'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [2:0] _exceptionNO_T_1 = io_memoryUnit_in_ex_exception_7 ? 3'h7 : _exceptionNO_T; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_2 = io_memoryUnit_in_ex_exception_13 ? 4'hd : {{1'd0}, _exceptionNO_T_1}; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_3 = io_memoryUnit_in_ex_exception_15 ? 4'hf : _exceptionNO_T_2; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_4 = io_memoryUnit_in_ex_exception_4 ? 4'h4 : _exceptionNO_T_3; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_5 = io_memoryUnit_in_ex_exception_6 ? 4'h6 : _exceptionNO_T_4; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_6 = io_memoryUnit_in_ex_exception_8 ? 4'h8 : _exceptionNO_T_5; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_7 = io_memoryUnit_in_ex_exception_9 ? 4'h9 : _exceptionNO_T_6; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_8 = io_memoryUnit_in_ex_exception_11 ? 4'hb : _exceptionNO_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_9 = io_memoryUnit_in_ex_exception_0 ? 4'h0 : _exceptionNO_T_8; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_10 = io_memoryUnit_in_ex_exception_2 ? 4'h2 : _exceptionNO_T_9; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_11 = io_memoryUnit_in_ex_exception_1 ? 4'h1 : _exceptionNO_T_10; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] _exceptionNO_T_12 = io_memoryUnit_in_ex_exception_12 ? 4'hc : _exceptionNO_T_11; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [3:0] exceptionNO = io_memoryUnit_in_ex_exception_3 ? 4'h3 : _exceptionNO_T_12; // @[playground/src/pipeline/execute/fu/Csr.scala 316:74]
  wire [2:0] _interruptNO_T = io_memoryUnit_in_ex_interrupt_4 ? 3'h4 : 3'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_1 = io_memoryUnit_in_ex_interrupt_8 ? 4'h8 : {{1'd0}, _interruptNO_T}; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_2 = io_memoryUnit_in_ex_interrupt_0 ? 4'h0 : _interruptNO_T_1; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_3 = io_memoryUnit_in_ex_interrupt_5 ? 4'h5 : _interruptNO_T_2; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_4 = io_memoryUnit_in_ex_interrupt_9 ? 4'h9 : _interruptNO_T_3; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_5 = io_memoryUnit_in_ex_interrupt_1 ? 4'h1 : _interruptNO_T_4; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_6 = io_memoryUnit_in_ex_interrupt_7 ? 4'h7 : _interruptNO_T_5; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] _interruptNO_T_7 = io_memoryUnit_in_ex_interrupt_11 ? 4'hb : _interruptNO_T_6; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [3:0] interruptNO = io_memoryUnit_in_ex_interrupt_3 ? 4'h3 : _interruptNO_T_7; // @[playground/src/pipeline/execute/fu/Csr.scala 317:74]
  wire [63:0] _causeNO_T = {raise_interrupt, 63'h0}; // @[playground/src/pipeline/execute/fu/Csr.scala 318:38]
  wire [3:0] _causeNO_T_1 = raise_interrupt ? interruptNO : exceptionNO; // @[playground/src/pipeline/execute/fu/Csr.scala 318:58]
  wire [63:0] _GEN_79 = {{60'd0}, _causeNO_T_1}; // @[playground/src/pipeline/execute/fu/Csr.scala 318:53]
  wire [63:0] causeNO = _causeNO_T | _GEN_79; // @[playground/src/pipeline/execute/fu/Csr.scala 318:53]
  wire [63:0] deleg = raise_interrupt ? mideleg : medeleg; // @[playground/src/pipeline/execute/fu/Csr.scala 320:19]
  wire [63:0] _delegS_T_1 = deleg >> causeNO[3:0]; // @[playground/src/pipeline/execute/fu/Csr.scala 321:22]
  wire  delegS = _delegS_T_1[0] & _interrupt_enable_0_T_6; // @[playground/src/pipeline/execute/fu/Csr.scala 321:59]
  wire  _tval_wen_T = ~raise_exception; // @[playground/src/pipeline/execute/fu/Csr.scala 324:5]
  wire  tval_wen = raise_interrupt | _tval_wen_T; // @[playground/src/pipeline/execute/fu/Csr.scala 323:34]
  wire [63:0] _GEN_25 = 4'h1 == exceptionNO ? io_memoryUnit_in_ex_tval_1 : io_memoryUnit_in_ex_tval_0; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_26 = 4'h2 == exceptionNO ? io_memoryUnit_in_ex_tval_2 : _GEN_25; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_27 = 4'h3 == exceptionNO ? io_memoryUnit_in_ex_tval_3 : _GEN_26; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_28 = 4'h4 == exceptionNO ? io_memoryUnit_in_ex_tval_4 : _GEN_27; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_29 = 4'h5 == exceptionNO ? io_memoryUnit_in_ex_tval_5 : _GEN_28; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_30 = 4'h6 == exceptionNO ? io_memoryUnit_in_ex_tval_6 : _GEN_29; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_31 = 4'h7 == exceptionNO ? io_memoryUnit_in_ex_tval_7 : _GEN_30; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_32 = 4'h8 == exceptionNO ? io_memoryUnit_in_ex_tval_8 : _GEN_31; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_33 = 4'h9 == exceptionNO ? io_memoryUnit_in_ex_tval_9 : _GEN_32; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_34 = 4'ha == exceptionNO ? io_memoryUnit_in_ex_tval_10 : _GEN_33; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_35 = 4'hb == exceptionNO ? io_memoryUnit_in_ex_tval_11 : _GEN_34; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_36 = 4'hc == exceptionNO ? io_memoryUnit_in_ex_tval_12 : _GEN_35; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_37 = 4'hd == exceptionNO ? io_memoryUnit_in_ex_tval_13 : _GEN_36; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_38 = 4'he == exceptionNO ? io_memoryUnit_in_ex_tval_14 : _GEN_37; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_39 = 4'hf == exceptionNO ? io_memoryUnit_in_ex_tval_15 : _GEN_38; // @[playground/src/pipeline/execute/fu/Csr.scala 329:{13,13}]
  wire [63:0] _GEN_40 = delegS ? _GEN_39 : _GEN_18; // @[playground/src/pipeline/execute/fu/Csr.scala 328:18 329:13]
  wire [63:0] _GEN_41 = delegS ? _GEN_20 : _GEN_39; // @[playground/src/pipeline/execute/fu/Csr.scala 328:18 331:13]
  wire [63:0] _GEN_42 = raise_exception ? _GEN_40 : _GEN_18; // @[playground/src/pipeline/execute/fu/Csr.scala 326:25]
  wire [63:0] _GEN_43 = raise_exception ? _GEN_41 : _GEN_20; // @[playground/src/pipeline/execute/fu/Csr.scala 326:25]
  wire [1:0] _GEN_48 = delegS ? mode : {{1'd0}, mstatusBundle_spp}; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 342:24 337:30]
  wire  mstatusNew_pie_s = delegS ? mstatusBundle_ie_s : mstatusBundle_pie_s; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 343:24 337:30]
  wire  mstatusNew_ie_s = delegS ? 1'h0 : mstatusBundle_ie_s; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 344:24 337:30]
  wire [1:0] _GEN_51 = delegS ? 2'h1 : 2'h3; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 345:24 353:24]
  wire [1:0] mstatusNew_mpp = delegS ? mstatusBundle_mpp : mode; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 337:30 350:24]
  wire  mstatusNew_pie_m = delegS ? mstatusBundle_pie_m : mstatusBundle_ie_m; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 337:30 351:24]
  wire  mstatusNew_ie_m = delegS & mstatusBundle_ie_m; // @[playground/src/pipeline/execute/fu/Csr.scala 339:18 337:30 352:24]
  wire [5:0] mstatus_lo_lo_1 = {mstatusNew_pie_s,mstatusBundle_pie_u,mstatusNew_ie_m,mstatusBundle_ie_h,mstatusNew_ie_s,
    mstatusBundle_ie_u}; // @[playground/src/pipeline/execute/fu/Csr.scala 356:27]
  wire  mstatusNew_spp = _GEN_48[0]; // @[playground/src/pipeline/execute/fu/Csr.scala 337:30]
  wire [14:0] mstatus_lo_1 = {mstatusBundle_fs,mstatusNew_mpp,mstatusBundle_hpp,mstatusNew_spp,mstatusNew_pie_m,
    mstatusBundle_pie_h,mstatus_lo_lo_1}; // @[playground/src/pipeline/execute/fu/Csr.scala 356:27]
  wire [6:0] mstatus_hi_lo_1 = {mstatusBundle_tw,mstatusBundle_tvm,mstatusBundle_mxr,mstatusBundle_sum,
    mstatusBundle_mprv,mstatusBundle_xs}; // @[playground/src/pipeline/execute/fu/Csr.scala 356:27]
  wire [63:0] _mstatus_T_9 = {mstatusBundle_sd,mstatusBundle_pad1,mstatusBundle_sxl,mstatusBundle_uxl,mstatusBundle_pad0
    ,mstatusBundle_tsr,mstatus_hi_lo_1,mstatus_lo_1}; // @[playground/src/pipeline/execute/fu/Csr.scala 356:27]
  wire [63:0] tvec = delegS ? stvec : mtvec; // @[playground/src/pipeline/execute/fu/Csr.scala 363:24]
  wire [63:0] _trap_target_T_1 = {tvec[63:2], 2'h0}; // @[playground/src/pipeline/execute/fu/Csr.scala 364:37]
  wire  _trap_target_T_3 = tvec[0] & raise_interrupt; // @[playground/src/pipeline/execute/fu/Csr.scala 365:13]
  wire [65:0] _trap_target_T_4 = {causeNO, 2'h0}; // @[playground/src/pipeline/execute/fu/Csr.scala 366:14]
  wire [65:0] _trap_target_T_5 = _trap_target_T_3 ? _trap_target_T_4 : 66'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 364:48]
  wire [65:0] _GEN_80 = {{2'd0}, _trap_target_T_1}; // @[playground/src/pipeline/execute/fu/Csr.scala 364:43]
  wire [65:0] _trap_target_T_7 = _GEN_80 + _trap_target_T_5; // @[playground/src/pipeline/execute/fu/Csr.scala 364:43]
  wire  mstatusNew_1_mprv = mstatusBundle_mpp != 2'h3 ? 1'h0 : mstatusBundle_mprv; // @[playground/src/pipeline/execute/fu/Csr.scala 373:36 374:23 372:30]
  wire [5:0] mstatus_lo_lo_2 = {mstatusBundle_pie_s,mstatusBundle_pie_u,mstatusBundle_pie_m,mstatusBundle_ie_h,
    mstatusBundle_ie_s,mstatusBundle_ie_u}; // @[playground/src/pipeline/execute/fu/Csr.scala 380:36]
  wire [14:0] mstatus_lo_2 = {mstatusBundle_fs,2'h0,mstatusBundle_hpp,mstatusBundle_spp,1'h1,mstatusBundle_pie_h,
    mstatus_lo_lo_2}; // @[playground/src/pipeline/execute/fu/Csr.scala 380:36]
  wire [6:0] mstatus_hi_lo_2 = {mstatusBundle_tw,mstatusBundle_tvm,mstatusBundle_mxr,mstatusBundle_sum,mstatusNew_1_mprv
    ,mstatusBundle_xs}; // @[playground/src/pipeline/execute/fu/Csr.scala 380:36]
  wire [63:0] _mstatus_T_10 = {mstatusBundle_sd,mstatusBundle_pad1,mstatusBundle_sxl,mstatusBundle_uxl,
    mstatusBundle_pad0,mstatusBundle_tsr,mstatus_hi_lo_2,mstatus_lo_2}; // @[playground/src/pipeline/execute/fu/Csr.scala 380:36]
  wire [1:0] _GEN_81 = {{1'd0}, mstatusBundle_spp}; // @[playground/src/pipeline/execute/fu/Csr.scala 388:25]
  wire  mstatusNew_2_mprv = _GEN_81 != 2'h3 ? 1'h0 : mstatusBundle_mprv; // @[playground/src/pipeline/execute/fu/Csr.scala 388:36 389:23 387:30]
  wire [1:0] _mode_T = {1'h0,mstatusBundle_spp}; // @[playground/src/pipeline/execute/fu/Csr.scala 392:28]
  wire [5:0] mstatus_lo_lo_3 = {1'h1,mstatusBundle_pie_u,mstatusBundle_ie_m,mstatusBundle_ie_h,mstatusBundle_pie_s,
    mstatusBundle_ie_u}; // @[playground/src/pipeline/execute/fu/Csr.scala 395:36]
  wire [14:0] mstatus_lo_3 = {mstatusBundle_fs,mstatusBundle_mpp,mstatusBundle_hpp,1'h0,mstatusBundle_pie_m,
    mstatusBundle_pie_h,mstatus_lo_lo_3}; // @[playground/src/pipeline/execute/fu/Csr.scala 395:36]
  wire [6:0] mstatus_hi_lo_3 = {mstatusBundle_tw,mstatusBundle_tvm,mstatusBundle_mxr,mstatusBundle_sum,mstatusNew_2_mprv
    ,mstatusBundle_xs}; // @[playground/src/pipeline/execute/fu/Csr.scala 395:36]
  wire [63:0] _mstatus_T_11 = {mstatusBundle_sd,mstatusBundle_pad1,mstatusBundle_sxl,mstatusBundle_uxl,
    mstatusBundle_pad0,mstatusBundle_tsr,mstatus_hi_lo_3,mstatus_lo_3}; // @[playground/src/pipeline/execute/fu/Csr.scala 395:36]
  wire [63:0] ret_target = isSret ? sepc : mepc; // @[playground/src/pipeline/execute/fu/Csr.scala 385:16 397:22]
  wire [63:0] trap_target = _trap_target_T_7[63:0]; // @[playground/src/pipeline/execute/fu/Csr.scala 362:25 364:15]
  assign io_decodeUnit_mode = mode; // @[playground/src/pipeline/execute/fu/Csr.scala 404:25]
  assign io_decodeUnit_interrupt = _io_decodeUnit_interrupt_T_2 & _io_decodeUnit_interrupt_T_3; // @[playground/src/pipeline/execute/fu/Csr.scala 258:79]
  assign io_executeUnit_out_rdata = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_executeUnit_out_ex_exception_1 = io_executeUnit_in_ex_exception_1; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_exception_2 = (illegal_addr | illegal_access) & write | io_executeUnit_in_ex_exception_2; // @[playground/src/pipeline/execute/fu/Csr.scala 407:47]
  assign io_executeUnit_out_ex_exception_3 = io_executeUnit_in_ex_exception_3; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_exception_8 = io_executeUnit_in_ex_exception_8; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_exception_9 = io_executeUnit_in_ex_exception_9; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_exception_11 = io_executeUnit_in_ex_exception_11; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_exception_12 = io_executeUnit_in_ex_exception_12; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_0 = io_executeUnit_in_ex_interrupt_0; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_1 = io_executeUnit_in_ex_interrupt_1; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_2 = io_executeUnit_in_ex_interrupt_2; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_3 = io_executeUnit_in_ex_interrupt_3; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_4 = io_executeUnit_in_ex_interrupt_4; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_5 = io_executeUnit_in_ex_interrupt_5; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_6 = io_executeUnit_in_ex_interrupt_6; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_7 = io_executeUnit_in_ex_interrupt_7; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_8 = io_executeUnit_in_ex_interrupt_8; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_9 = io_executeUnit_in_ex_interrupt_9; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_10 = io_executeUnit_in_ex_interrupt_10; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_interrupt_11 = io_executeUnit_in_ex_interrupt_11; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_tval_1 = io_executeUnit_in_ex_tval_1; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_ex_tval_2 = io_executeUnit_in_info_inst; // @[playground/src/pipeline/execute/fu/Csr.scala 408:43]
  assign io_executeUnit_out_ex_tval_12 = io_executeUnit_in_ex_tval_12; // @[playground/src/pipeline/execute/fu/Csr.scala 405:25]
  assign io_executeUnit_out_flush = _T_105 & write; // @[playground/src/pipeline/execute/fu/Csr.scala 302:40]
  assign io_executeUnit_out_target = io_executeUnit_in_pc + 64'h4; // @[playground/src/pipeline/execute/fu/Csr.scala 411:68]
  assign io_memoryUnit_out_flush = raise_exc_int | ret; // @[playground/src/pipeline/execute/fu/Csr.scala 412:61]
  assign io_memoryUnit_out_target = raise_exc_int ? trap_target : ret_target; // @[playground/src/pipeline/execute/fu/Csr.scala 413:50]
  assign io_memoryUnit_out_lr = lr; // @[playground/src/pipeline/execute/fu/Csr.scala 162:29]
  assign io_memoryUnit_out_lr_addr = lr_addr; // @[playground/src/pipeline/execute/fu/Csr.scala 163:29]
  assign io_tlb_satp = satp; // @[playground/src/pipeline/execute/fu/Csr.scala 402:25]
  assign io_tlb_mstatus = mstatus; // @[playground/src/pipeline/execute/fu/Csr.scala 403:25]
  assign io_tlb_imode = mode; // @[playground/src/pipeline/execute/fu/Csr.scala 400:25]
  assign io_tlb_dmode = mstatusBundle_mprv ? mstatusBundle_mpp : mode; // @[playground/src/pipeline/execute/fu/Csr.scala 401:31]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 81:26]
      mstatus <= 64'ha00000000; // @[playground/src/pipeline/execute/fu/Csr.scala 81:26]
    end else if (isSret) begin // @[playground/src/pipeline/execute/fu/Csr.scala 385:16]
      mstatus <= _mstatus_T_11; // @[playground/src/pipeline/execute/fu/Csr.scala 395:22]
    end else if (isMret) begin // @[playground/src/pipeline/execute/fu/Csr.scala 370:16]
      mstatus <= _mstatus_T_10; // @[playground/src/pipeline/execute/fu/Csr.scala 380:22]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      mstatus <= _mstatus_T_9; // @[playground/src/pipeline/execute/fu/Csr.scala 356:13]
    end else begin
      mstatus <= _GEN_9;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 93:27]
      medeleg <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 93:27]
    end else if (wen & addr == 12'h302) begin // @[playground/src/defines/Util.scala 115:73]
      medeleg <= _medeleg_T_3; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 94:27]
      mideleg <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 94:27]
    end else if (wen & addr == 12'h303) begin // @[playground/src/defines/Util.scala 115:73]
      mideleg <= _mideleg_T_3; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 95:27]
      mie <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 95:27]
    end else if (wen & addr == 12'h304) begin // @[playground/src/defines/Util.scala 115:73]
      mie <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end else if (wen & addr == 12'h104) begin // @[playground/src/defines/Util.scala 115:73]
      mie <= _mie_T_3; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 96:27]
      mtvec <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 96:27]
    end else if (wen & addr == 12'h305) begin // @[playground/src/defines/Util.scala 115:73]
      mtvec <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 97:27]
      mcounteren <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 97:27]
    end else if (wen & addr == 12'h306) begin // @[playground/src/defines/Util.scala 115:73]
      mcounteren <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 100:27]
      mscratch <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 100:27]
    end else if (wen & addr == 12'h340) begin // @[playground/src/defines/Util.scala 115:73]
      mscratch <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 101:27]
      mepc <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 101:27]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      if (delegS) begin // @[playground/src/pipeline/execute/fu/Csr.scala 339:18]
        mepc <= _GEN_19;
      end else begin
        mepc <= io_memoryUnit_in_pc; // @[playground/src/pipeline/execute/fu/Csr.scala 349:24]
      end
    end else begin
      mepc <= _GEN_19;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 102:27]
      mcause <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 102:27]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      if (delegS) begin // @[playground/src/pipeline/execute/fu/Csr.scala 339:18]
        mcause <= _GEN_17;
      end else begin
        mcause <= causeNO; // @[playground/src/pipeline/execute/fu/Csr.scala 348:24]
      end
    end else begin
      mcause <= _GEN_17;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 103:27]
      mtval <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 103:27]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      if (delegS) begin // @[playground/src/pipeline/execute/fu/Csr.scala 339:18]
        mtval <= _GEN_43;
      end else if (tval_wen) begin // @[playground/src/pipeline/execute/fu/Csr.scala 354:22]
        mtval <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 354:30]
      end else begin
        mtval <= _GEN_43;
      end
    end else begin
      mtval <= _GEN_43;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 105:27]
      mipReg <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 105:27]
    end else if (wen & addr == 12'h144) begin // @[playground/src/defines/Util.scala 115:73]
      mipReg <= _mipReg_T_7; // @[playground/src/defines/Util.scala 115:77]
    end else if (wen & addr == 12'h344) begin // @[playground/src/defines/Util.scala 115:73]
      mipReg <= _mipReg_T_3; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 122:23]
      mcycle <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 122:23]
    end else if (wen & addr == 12'hc00) begin // @[playground/src/defines/Util.scala 115:73]
      mcycle <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end else begin
      mcycle <= _mcycle_T_1; // @[playground/src/pipeline/execute/fu/Csr.scala 123:10]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 134:27]
      stvec <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 134:27]
    end else if (wen & addr == 12'h105) begin // @[playground/src/defines/Util.scala 115:73]
      stvec <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 135:27]
      scounteren <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 135:27]
    end else if (wen & addr == 12'h106) begin // @[playground/src/defines/Util.scala 115:73]
      scounteren <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 138:25]
      sscratch <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 138:25]
    end else if (wen & addr == 12'h140) begin // @[playground/src/defines/Util.scala 115:73]
      sscratch <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 139:25]
      sepc <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 139:25]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      if (delegS) begin // @[playground/src/pipeline/execute/fu/Csr.scala 339:18]
        sepc <= io_memoryUnit_in_pc; // @[playground/src/pipeline/execute/fu/Csr.scala 341:24]
      end else begin
        sepc <= _GEN_16;
      end
    end else begin
      sepc <= _GEN_16;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 140:25]
      scause <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 140:25]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      if (delegS) begin // @[playground/src/pipeline/execute/fu/Csr.scala 339:18]
        scause <= causeNO; // @[playground/src/pipeline/execute/fu/Csr.scala 340:24]
      end else begin
        scause <= _GEN_12;
      end
    end else begin
      scause <= _GEN_12;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 141:25]
      stval <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 141:25]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      if (delegS) begin // @[playground/src/pipeline/execute/fu/Csr.scala 339:18]
        if (tval_wen) begin // @[playground/src/pipeline/execute/fu/Csr.scala 346:22]
          stval <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 346:30]
        end else begin
          stval <= _GEN_42;
        end
      end else begin
        stval <= _GEN_42;
      end
    end else begin
      stval <= _GEN_42;
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 146:21]
      satp <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 146:21]
    end else if (wen & addr == 12'h180) begin // @[playground/src/defines/Util.scala 115:73]
      satp <= wdata; // @[playground/src/defines/Util.scala 115:77]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 159:25]
      lr <= 1'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 159:25]
    end else if (isSret) begin // @[playground/src/pipeline/execute/fu/Csr.scala 385:16]
      lr <= 1'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 396:22]
    end else if (isMret) begin // @[playground/src/pipeline/execute/fu/Csr.scala 370:16]
      lr <= 1'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 381:22]
    end else if (io_memoryUnit_in_lr_wen) begin // @[playground/src/pipeline/execute/fu/Csr.scala 165:16]
      lr <= io_memoryUnit_in_lr_wbit; // @[playground/src/pipeline/execute/fu/Csr.scala 166:13]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 160:25]
      lr_addr <= 64'h0; // @[playground/src/pipeline/execute/fu/Csr.scala 160:25]
    end else if (io_memoryUnit_in_lr_wen) begin // @[playground/src/pipeline/execute/fu/Csr.scala 165:16]
      lr_addr <= io_memoryUnit_in_lr_waddr; // @[playground/src/pipeline/execute/fu/Csr.scala 167:13]
    end
    if (reset) begin // @[playground/src/pipeline/execute/fu/Csr.scala 234:21]
      mode <= 2'h3; // @[playground/src/pipeline/execute/fu/Csr.scala 234:21]
    end else if (isSret) begin // @[playground/src/pipeline/execute/fu/Csr.scala 385:16]
      mode <= _mode_T; // @[playground/src/pipeline/execute/fu/Csr.scala 392:22]
    end else if (isMret) begin // @[playground/src/pipeline/execute/fu/Csr.scala 370:16]
      mode <= mstatusBundle_mpp; // @[playground/src/pipeline/execute/fu/Csr.scala 377:22]
    end else if (raise_exc_int) begin // @[playground/src/pipeline/execute/fu/Csr.scala 335:23]
      mode <= _GEN_51;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mstatus = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  medeleg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mideleg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mie = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtvec = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mcounteren = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mscratch = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mepc = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mcause = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  mtval = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mipReg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mcycle = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  stvec = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  scounteren = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  sscratch = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  sepc = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  scause = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  stval = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  satp = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  lr = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  lr_addr = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  mode = _RAND_21[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemoryStage(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_ctrl_clear, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_pc, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_info_valid, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [2:0]  io_executeUnit_inst_0_info_fusel, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [6:0]  io_executeUnit_inst_0_info_op, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_info_reg_wen, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [4:0]  io_executeUnit_inst_0_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_info_imm, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_info_inst, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_exception_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_0_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_ex_tval_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_ex_tval_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_ex_tval_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_0_ex_tval_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_pc, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_info_valid, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [2:0]  io_executeUnit_inst_1_info_fusel, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [6:0]  io_executeUnit_inst_1_info_op, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_info_reg_wen, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [4:0]  io_executeUnit_inst_1_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_info_imm, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_info_inst, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_exception_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input         io_executeUnit_inst_1_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_ex_tval_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_ex_tval_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_ex_tval_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  input  [63:0] io_executeUnit_inst_1_ex_tval_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_pc, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_info_valid, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [2:0]  io_memoryUnit_inst_0_info_fusel, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [6:0]  io_memoryUnit_inst_0_info_op, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_info_reg_wen, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [4:0]  io_memoryUnit_inst_0_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_info_imm, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_info_inst, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_exception_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_0_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_ex_tval_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_ex_tval_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_ex_tval_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_0_ex_tval_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_pc, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_info_valid, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [2:0]  io_memoryUnit_inst_1_info_fusel, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [6:0]  io_memoryUnit_inst_1_info_op, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_info_reg_wen, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [4:0]  io_memoryUnit_inst_1_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_info_imm, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_info_inst, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_exception_12, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output        io_memoryUnit_inst_1_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_ex_tval_0, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_ex_tval_1, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_ex_tval_2, // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
  output [63:0] io_memoryUnit_inst_1_ex_tval_12 // @[playground/src/pipeline/memory/MemoryStage.scala 22:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] inst_0_pc; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_info_valid; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [2:0] inst_0_info_fusel; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [6:0] inst_0_info_op; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_info_reg_wen; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [4:0] inst_0_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_info_imm; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_info_inst; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_1; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_3; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_8; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_9; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_11; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_exception_12; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_0_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_ex_tval_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_ex_tval_1; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_ex_tval_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_0_ex_tval_12; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_pc; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_info_valid; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [2:0] inst_1_info_fusel; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [6:0] inst_1_info_op; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_info_reg_wen; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [4:0] inst_1_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_info_imm; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_info_inst; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_1; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_3; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_8; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_9; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_11; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_exception_12; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg  inst_1_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_ex_tval_0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_ex_tval_1; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_ex_tval_2; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  reg [63:0] inst_1_ex_tval_12; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
  assign io_memoryUnit_inst_0_pc = inst_0_pc; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_valid = inst_0_info_valid; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_fusel = inst_0_info_fusel; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_op = inst_0_info_op; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_reg_wen = inst_0_info_reg_wen; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_reg_waddr = inst_0_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_imm = inst_0_info_imm; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_info_inst = inst_0_info_inst; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_rd_info_wdata_0 = inst_0_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_rd_info_wdata_2 = inst_0_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_rd_info_wdata_3 = inst_0_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_rd_info_wdata_5 = inst_0_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_src_info_src1_data = inst_0_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_src_info_src2_data = inst_0_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_0 = inst_0_ex_exception_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_1 = inst_0_ex_exception_1; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_2 = inst_0_ex_exception_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_3 = inst_0_ex_exception_3; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_8 = inst_0_ex_exception_8; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_9 = inst_0_ex_exception_9; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_11 = inst_0_ex_exception_11; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_exception_12 = inst_0_ex_exception_12; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_0 = inst_0_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_1 = inst_0_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_2 = inst_0_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_3 = inst_0_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_4 = inst_0_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_5 = inst_0_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_6 = inst_0_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_7 = inst_0_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_8 = inst_0_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_9 = inst_0_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_10 = inst_0_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_interrupt_11 = inst_0_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_tval_0 = inst_0_ex_tval_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_tval_1 = inst_0_ex_tval_1; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_tval_2 = inst_0_ex_tval_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_0_ex_tval_12 = inst_0_ex_tval_12; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_pc = inst_1_pc; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_valid = inst_1_info_valid; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_fusel = inst_1_info_fusel; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_op = inst_1_info_op; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_reg_wen = inst_1_info_reg_wen; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_reg_waddr = inst_1_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_imm = inst_1_info_imm; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_info_inst = inst_1_info_inst; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_rd_info_wdata_0 = inst_1_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_rd_info_wdata_2 = inst_1_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_rd_info_wdata_3 = inst_1_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_rd_info_wdata_5 = inst_1_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_src_info_src1_data = inst_1_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_src_info_src2_data = inst_1_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_0 = inst_1_ex_exception_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_1 = inst_1_ex_exception_1; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_2 = inst_1_ex_exception_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_3 = inst_1_ex_exception_3; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_8 = inst_1_ex_exception_8; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_9 = inst_1_ex_exception_9; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_11 = inst_1_ex_exception_11; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_exception_12 = inst_1_ex_exception_12; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_0 = inst_1_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_1 = inst_1_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_2 = inst_1_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_3 = inst_1_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_4 = inst_1_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_5 = inst_1_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_6 = inst_1_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_7 = inst_1_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_8 = inst_1_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_9 = inst_1_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_10 = inst_1_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_interrupt_11 = inst_1_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_tval_0 = inst_1_ex_tval_0; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_tval_1 = inst_1_ex_tval_1; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_tval_2 = inst_1_ex_tval_2; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  assign io_memoryUnit_inst_1_ex_tval_12 = inst_1_ex_tval_12; // @[playground/src/pipeline/memory/MemoryStage.scala 40:22]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_pc <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_pc <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_pc <= io_executeUnit_inst_0_pc; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_valid <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_valid <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_valid <= io_executeUnit_inst_0_info_valid; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_fusel <= 3'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_fusel <= 3'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_fusel <= io_executeUnit_inst_0_info_fusel; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_op <= 7'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_op <= 7'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_op <= io_executeUnit_inst_0_info_op; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_reg_wen <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_reg_wen <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_reg_wen <= io_executeUnit_inst_0_info_reg_wen; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_reg_waddr <= io_executeUnit_inst_0_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_imm <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_imm <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_imm <= io_executeUnit_inst_0_info_imm; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_info_inst <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_info_inst <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_info_inst <= io_executeUnit_inst_0_info_inst; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_rd_info_wdata_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_rd_info_wdata_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_rd_info_wdata_0 <= io_executeUnit_inst_0_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_rd_info_wdata_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_rd_info_wdata_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_rd_info_wdata_2 <= io_executeUnit_inst_0_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_rd_info_wdata_3 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_rd_info_wdata_3 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_rd_info_wdata_3 <= io_executeUnit_inst_0_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_rd_info_wdata_5 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_rd_info_wdata_5 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_rd_info_wdata_5 <= io_executeUnit_inst_0_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_src_info_src1_data <= io_executeUnit_inst_0_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_src_info_src2_data <= io_executeUnit_inst_0_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_0 <= io_executeUnit_inst_0_ex_exception_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_1 <= io_executeUnit_inst_0_ex_exception_1; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_2 <= io_executeUnit_inst_0_ex_exception_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_3 <= io_executeUnit_inst_0_ex_exception_3; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_8 <= io_executeUnit_inst_0_ex_exception_8; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_9 <= io_executeUnit_inst_0_ex_exception_9; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_11 <= io_executeUnit_inst_0_ex_exception_11; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_exception_12 <= io_executeUnit_inst_0_ex_exception_12; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_0 <= io_executeUnit_inst_0_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_1 <= io_executeUnit_inst_0_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_2 <= io_executeUnit_inst_0_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_3 <= io_executeUnit_inst_0_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_4 <= io_executeUnit_inst_0_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_5 <= io_executeUnit_inst_0_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_6 <= io_executeUnit_inst_0_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_7 <= io_executeUnit_inst_0_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_8 <= io_executeUnit_inst_0_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_9 <= io_executeUnit_inst_0_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_10 <= io_executeUnit_inst_0_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_interrupt_11 <= io_executeUnit_inst_0_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_tval_0 <= io_executeUnit_inst_0_ex_tval_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_tval_1 <= io_executeUnit_inst_0_ex_tval_1; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_tval_2 <= io_executeUnit_inst_0_ex_tval_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_0_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_0_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_0_ex_tval_12 <= io_executeUnit_inst_0_ex_tval_12; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_pc <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_pc <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_pc <= io_executeUnit_inst_1_pc; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_valid <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_valid <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_valid <= io_executeUnit_inst_1_info_valid; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_fusel <= 3'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_fusel <= 3'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_fusel <= io_executeUnit_inst_1_info_fusel; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_op <= 7'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_op <= 7'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_op <= io_executeUnit_inst_1_info_op; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_reg_wen <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_reg_wen <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_reg_wen <= io_executeUnit_inst_1_info_reg_wen; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_reg_waddr <= io_executeUnit_inst_1_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_imm <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_imm <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_imm <= io_executeUnit_inst_1_info_imm; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_info_inst <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_info_inst <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_info_inst <= io_executeUnit_inst_1_info_inst; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_rd_info_wdata_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_rd_info_wdata_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_rd_info_wdata_0 <= io_executeUnit_inst_1_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_rd_info_wdata_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_rd_info_wdata_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_rd_info_wdata_2 <= io_executeUnit_inst_1_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_rd_info_wdata_3 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_rd_info_wdata_3 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_rd_info_wdata_3 <= io_executeUnit_inst_1_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_rd_info_wdata_5 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_rd_info_wdata_5 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_rd_info_wdata_5 <= io_executeUnit_inst_1_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_src_info_src1_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_src_info_src1_data <= io_executeUnit_inst_1_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_src_info_src2_data <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_src_info_src2_data <= io_executeUnit_inst_1_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_0 <= io_executeUnit_inst_1_ex_exception_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_1 <= io_executeUnit_inst_1_ex_exception_1; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_2 <= io_executeUnit_inst_1_ex_exception_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_3 <= io_executeUnit_inst_1_ex_exception_3; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_8 <= io_executeUnit_inst_1_ex_exception_8; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_9 <= io_executeUnit_inst_1_ex_exception_9; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_11 <= io_executeUnit_inst_1_ex_exception_11; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_exception_12 <= io_executeUnit_inst_1_ex_exception_12; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_0 <= io_executeUnit_inst_1_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_1 <= io_executeUnit_inst_1_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_2 <= io_executeUnit_inst_1_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_3 <= io_executeUnit_inst_1_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_4 <= io_executeUnit_inst_1_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_5 <= io_executeUnit_inst_1_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_6 <= io_executeUnit_inst_1_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_7 <= io_executeUnit_inst_1_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_8 <= io_executeUnit_inst_1_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_9 <= io_executeUnit_inst_1_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_10 <= io_executeUnit_inst_1_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_interrupt_11 <= io_executeUnit_inst_1_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_tval_0 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_tval_0 <= io_executeUnit_inst_1_ex_tval_0; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_tval_1 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_tval_1 <= io_executeUnit_inst_1_ex_tval_1; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_tval_2 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_tval_2 <= io_executeUnit_inst_1_ex_tval_2; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
    if (reset) begin // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
      inst_1_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 30:51]
    end else if (io_ctrl_clear) begin // @[playground/src/pipeline/memory/MemoryStage.scala 33:25]
      inst_1_ex_tval_12 <= 64'h0; // @[playground/src/pipeline/memory/MemoryStage.scala 34:15]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/memory/MemoryStage.scala 35:37]
      inst_1_ex_tval_12 <= io_executeUnit_inst_1_ex_tval_12; // @[playground/src/pipeline/memory/MemoryStage.scala 36:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  inst_0_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  inst_0_info_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_0_info_fusel = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  inst_0_info_op = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  inst_0_info_reg_wen = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  inst_0_info_reg_waddr = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  inst_0_info_imm = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  inst_0_info_inst = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  inst_0_rd_info_wdata_0 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  inst_0_rd_info_wdata_2 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  inst_0_rd_info_wdata_3 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  inst_0_rd_info_wdata_5 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  inst_0_src_info_src1_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  inst_0_src_info_src2_data = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  inst_0_ex_exception_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inst_0_ex_exception_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  inst_0_ex_exception_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  inst_0_ex_exception_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  inst_0_ex_exception_8 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  inst_0_ex_exception_9 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inst_0_ex_exception_11 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  inst_0_ex_exception_12 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  inst_0_ex_interrupt_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  inst_0_ex_interrupt_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  inst_0_ex_interrupt_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  inst_0_ex_interrupt_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  inst_0_ex_interrupt_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  inst_0_ex_interrupt_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  inst_0_ex_interrupt_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inst_0_ex_interrupt_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  inst_0_ex_interrupt_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  inst_0_ex_interrupt_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  inst_0_ex_interrupt_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  inst_0_ex_interrupt_11 = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  inst_0_ex_tval_0 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  inst_0_ex_tval_1 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  inst_0_ex_tval_2 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  inst_0_ex_tval_12 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  inst_1_pc = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  inst_1_info_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  inst_1_info_fusel = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  inst_1_info_op = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  inst_1_info_reg_wen = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  inst_1_info_reg_waddr = _RAND_43[4:0];
  _RAND_44 = {2{`RANDOM}};
  inst_1_info_imm = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  inst_1_info_inst = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  inst_1_rd_info_wdata_0 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  inst_1_rd_info_wdata_2 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  inst_1_rd_info_wdata_3 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  inst_1_rd_info_wdata_5 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  inst_1_src_info_src1_data = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  inst_1_src_info_src2_data = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  inst_1_ex_exception_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  inst_1_ex_exception_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  inst_1_ex_exception_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  inst_1_ex_exception_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  inst_1_ex_exception_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  inst_1_ex_exception_9 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  inst_1_ex_exception_11 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  inst_1_ex_exception_12 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  inst_1_ex_interrupt_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  inst_1_ex_interrupt_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  inst_1_ex_interrupt_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  inst_1_ex_interrupt_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  inst_1_ex_interrupt_4 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  inst_1_ex_interrupt_5 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  inst_1_ex_interrupt_6 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  inst_1_ex_interrupt_7 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  inst_1_ex_interrupt_8 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  inst_1_ex_interrupt_9 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  inst_1_ex_interrupt_10 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  inst_1_ex_interrupt_11 = _RAND_71[0:0];
  _RAND_72 = {2{`RANDOM}};
  inst_1_ex_tval_0 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  inst_1_ex_tval_1 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  inst_1_ex_tval_2 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  inst_1_ex_tval_12 = _RAND_75[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AtomAlu(
  input  [63:0] io_in_rdata, // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 10:14]
  input  [63:0] io_in_src2, // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 10:14]
  input  [6:0]  io_in_info_op, // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 10:14]
  input  [63:0] io_in_info_inst, // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 10:14]
  output [63:0] io_out_result // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 10:14]
);
  wire  is_sub = ~io_in_info_op[6]; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 24:17]
  wire [63:0] _sum_T_1 = is_sub ? 64'hffffffffffffffff : 64'h0; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 25:38]
  wire [63:0] _sum_T_2 = io_in_src2 ^ _sum_T_1; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 25:32]
  wire [64:0] _sum_T_3 = io_in_rdata + _sum_T_2; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 25:23]
  wire [64:0] _GEN_0 = {{64'd0}, is_sub}; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 25:55]
  wire [64:0] sum = _sum_T_3 + _GEN_0; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 25:55]
  wire [63:0] oxr = io_in_rdata ^ io_in_src2; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 26:22]
  wire  sltu = ~sum[64]; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 27:17]
  wire  slt = oxr[63] ^ sltu; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 28:31]
  wire  is_word = ~io_in_info_inst[12]; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 29:17]
  wire [63:0] _res_T_1 = io_in_rdata & io_in_src2; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 38:34]
  wire [63:0] _res_T_2 = io_in_rdata | io_in_src2; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 39:34]
  wire [63:0] _res_T_4 = slt ? io_in_rdata : io_in_src2; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 40:31]
  wire [63:0] _res_T_6 = slt ? io_in_src2 : io_in_rdata; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 41:31]
  wire [63:0] _res_T_8 = sltu ? io_in_rdata : io_in_src2; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 42:31]
  wire [63:0] _res_T_10 = sltu ? io_in_src2 : io_in_rdata; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 43:31]
  wire [64:0] _res_T_12 = 6'h22 == io_in_info_op[5:0] ? {{1'd0}, io_in_src2} : sum; // @[playground/src/defines/Util.scala 51:28]
  wire [6:0] _GEN_1 = {{1'd0}, io_in_info_op[5:0]}; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_14 = 7'h63 == _GEN_1 ? sum : _res_T_12; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_16 = 6'h24 == io_in_info_op[5:0] ? {{1'd0}, oxr} : _res_T_14; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_18 = 6'h25 == io_in_info_op[5:0] ? {{1'd0}, _res_T_1} : _res_T_16; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_20 = 6'h26 == io_in_info_op[5:0] ? {{1'd0}, _res_T_2} : _res_T_18; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_22 = 6'h37 == io_in_info_op[5:0] ? {{1'd0}, _res_T_4} : _res_T_20; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_24 = 6'h30 == io_in_info_op[5:0] ? {{1'd0}, _res_T_6} : _res_T_22; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] _res_T_26 = 6'h31 == io_in_info_op[5:0] ? {{1'd0}, _res_T_8} : _res_T_24; // @[playground/src/defines/Util.scala 51:28]
  wire [64:0] res = 6'h32 == io_in_info_op[5:0] ? {{1'd0}, _res_T_10} : _res_T_26; // @[playground/src/defines/Util.scala 51:28]
  wire  io_out_result_signBit = res[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _io_out_result_T_2 = io_out_result_signBit ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _io_out_result_T_3 = {_io_out_result_T_2,res[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  assign io_out_result = is_word ? _io_out_result_T_3 : res[63:0]; // @[playground/src/pipeline/memory/lsu/AtomAlu.scala 47:23]
endmodule
module LsExecute(
  input         io_dataMemory_in_access_fault, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input         io_dataMemory_in_page_fault, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input         io_dataMemory_in_ready, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input  [63:0] io_dataMemory_in_rdata, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output        io_dataMemory_out_en, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output [7:0]  io_dataMemory_out_rlen, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output        io_dataMemory_out_wen, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output [7:0]  io_dataMemory_out_wstrb, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output [63:0] io_dataMemory_out_addr, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output [63:0] io_dataMemory_out_wdata, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input         io_in_mem_en, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input  [63:0] io_in_mem_addr, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input  [63:0] io_in_wdata, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  input  [6:0]  io_in_info_op, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output        io_out_addr_misaligned, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output        io_out_access_fault, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output        io_out_page_fault, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output [63:0] io_out_rdata, // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
  output        io_out_ready // @[playground/src/pipeline/memory/lsu/LsExecute.scala 10:14]
);
  wire  is_store = io_in_mem_en & io_in_info_op[3]; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 75:28]
  wire  partial_load = ~is_store & io_in_info_op != 7'h3; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 76:32]
  wire [1:0] size = io_in_info_op[1:0]; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 78:21]
  wire [63:0] _req_wdata_T_3 = {io_in_wdata[7:0],io_in_wdata[7:0],io_in_wdata[7:0],io_in_wdata[7:0],io_in_wdata[7:0],
    io_in_wdata[7:0],io_in_wdata[7:0],io_in_wdata[7:0]}; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 42:24]
  wire [63:0] _req_wdata_T_6 = {io_in_wdata[15:0],io_in_wdata[15:0],io_in_wdata[15:0],io_in_wdata[15:0]}; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 43:24]
  wire [63:0] _req_wdata_T_8 = {io_in_wdata[31:0],io_in_wdata[31:0]}; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 44:24]
  wire  _req_wdata_T_9 = 2'h0 == size; // @[playground/src/defines/Util.scala 46:34]
  wire  _req_wdata_T_10 = 2'h1 == size; // @[playground/src/defines/Util.scala 46:34]
  wire  _req_wdata_T_11 = 2'h2 == size; // @[playground/src/defines/Util.scala 46:34]
  wire  _req_wdata_T_12 = 2'h3 == size; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _req_wdata_T_13 = _req_wdata_T_9 ? _req_wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _req_wdata_T_14 = _req_wdata_T_10 ? _req_wdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _req_wdata_T_15 = _req_wdata_T_11 ? _req_wdata_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _req_wdata_T_16 = _req_wdata_T_12 ? io_in_wdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _req_wdata_T_17 = _req_wdata_T_13 | _req_wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _req_wdata_T_18 = _req_wdata_T_17 | _req_wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _req_wmask_T_5 = _req_wdata_T_10 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _req_wmask_T_6 = _req_wdata_T_11 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _req_wmask_T_7 = _req_wdata_T_12 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_0 = {{1'd0}, _req_wdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _req_wmask_T_8 = _GEN_0 | _req_wmask_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _GEN_1 = {{2'd0}, _req_wmask_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _req_wmask_T_9 = _GEN_1 | _req_wmask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _GEN_2 = {{4'd0}, _req_wmask_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _req_wmask_T_10 = _GEN_2 | _req_wmask_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [14:0] _GEN_10 = {{7'd0}, _req_wmask_T_10}; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 36:7]
  wire [14:0] req_wmask = _GEN_10 << io_in_mem_addr[2:0]; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 36:7]
  wire  _rdata64_T_9 = 3'h0 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_10 = 3'h1 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_11 = 3'h2 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_12 = 3'h3 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_13 = 3'h4 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_14 = 3'h5 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_15 = 3'h6 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata64_T_16 = 3'h7 == io_in_mem_addr[2:0]; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata64_T_17 = _rdata64_T_9 ? io_dataMemory_in_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [55:0] _rdata64_T_18 = _rdata64_T_10 ? io_dataMemory_in_rdata[63:8] : 56'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [47:0] _rdata64_T_19 = _rdata64_T_11 ? io_dataMemory_in_rdata[63:16] : 48'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [39:0] _rdata64_T_20 = _rdata64_T_12 ? io_dataMemory_in_rdata[63:24] : 40'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata64_T_21 = _rdata64_T_13 ? io_dataMemory_in_rdata[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [23:0] _rdata64_T_22 = _rdata64_T_14 ? io_dataMemory_in_rdata[63:40] : 24'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _rdata64_T_23 = _rdata64_T_15 ? io_dataMemory_in_rdata[63:48] : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdata64_T_24 = _rdata64_T_16 ? io_dataMemory_in_rdata[63:56] : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_3 = {{8'd0}, _rdata64_T_18}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata64_T_25 = _rdata64_T_17 | _GEN_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_4 = {{16'd0}, _rdata64_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata64_T_26 = _rdata64_T_25 | _GEN_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_5 = {{24'd0}, _rdata64_T_20}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata64_T_27 = _rdata64_T_26 | _GEN_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_6 = {{32'd0}, _rdata64_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata64_T_28 = _rdata64_T_27 | _GEN_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_7 = {{40'd0}, _rdata64_T_22}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata64_T_29 = _rdata64_T_28 | _GEN_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_8 = {{48'd0}, _rdata64_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata64_T_30 = _rdata64_T_29 | _GEN_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_9 = {{56'd0}, _rdata64_T_24}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata64 = _rdata64_T_30 | _GEN_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  rdata_partial_result_signBit = rdata64[7]; // @[playground/src/defines/Util.scala 33:20]
  wire [55:0] _rdata_partial_result_T_2 = rdata_partial_result_signBit ? 56'hffffffffffffff : 56'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _rdata_partial_result_T_3 = {_rdata_partial_result_T_2,rdata64[7:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire  rdata_partial_result_signBit_1 = rdata64[15]; // @[playground/src/defines/Util.scala 33:20]
  wire [47:0] _rdata_partial_result_T_6 = rdata_partial_result_signBit_1 ? 48'hffffffffffff : 48'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _rdata_partial_result_T_7 = {_rdata_partial_result_T_6,rdata64[15:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire  rdata_partial_result_signBit_2 = rdata64[31]; // @[playground/src/defines/Util.scala 33:20]
  wire [31:0] _rdata_partial_result_T_10 = rdata_partial_result_signBit_2 ? 32'hffffffff : 32'h0; // @[playground/src/defines/Util.scala 34:49]
  wire [63:0] _rdata_partial_result_T_11 = {_rdata_partial_result_T_10,rdata64[31:0]}; // @[playground/src/defines/Util.scala 34:44]
  wire [63:0] _rdata_partial_result_T_13 = {56'h0,rdata64[7:0]}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _rdata_partial_result_T_15 = {48'h0,rdata64[15:0]}; // @[playground/src/defines/Util.scala 41:44]
  wire [63:0] _rdata_partial_result_T_17 = {32'h0,rdata64[31:0]}; // @[playground/src/defines/Util.scala 41:44]
  wire  _rdata_partial_result_T_18 = 7'h0 == io_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_partial_result_T_19 = 7'h1 == io_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_partial_result_T_20 = 7'h2 == io_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_partial_result_T_21 = 7'h4 == io_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_partial_result_T_22 = 7'h5 == io_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire  _rdata_partial_result_T_23 = 7'h6 == io_in_info_op; // @[playground/src/defines/Util.scala 46:34]
  wire [63:0] _rdata_partial_result_T_24 = _rdata_partial_result_T_18 ? _rdata_partial_result_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_25 = _rdata_partial_result_T_19 ? _rdata_partial_result_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_26 = _rdata_partial_result_T_20 ? _rdata_partial_result_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_27 = _rdata_partial_result_T_21 ? _rdata_partial_result_T_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_28 = _rdata_partial_result_T_22 ? _rdata_partial_result_T_15 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_29 = _rdata_partial_result_T_23 ? _rdata_partial_result_T_17 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_30 = _rdata_partial_result_T_24 | _rdata_partial_result_T_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_31 = _rdata_partial_result_T_30 | _rdata_partial_result_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_32 = _rdata_partial_result_T_31 | _rdata_partial_result_T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_partial_result_T_33 = _rdata_partial_result_T_32 | _rdata_partial_result_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata_partial_result = _rdata_partial_result_T_33 | _rdata_partial_result_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _addr_aligned_T_2 = ~io_in_mem_addr[0]; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 125:27]
  wire  _addr_aligned_T_4 = io_in_mem_addr[1:0] == 2'h0; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 126:30]
  wire  _addr_aligned_T_6 = io_in_mem_addr[2:0] == 3'h0; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 127:30]
  wire  addr_aligned = _req_wdata_T_9 | _req_wdata_T_10 & _addr_aligned_T_2 | _req_wdata_T_11 & _addr_aligned_T_4 |
    _req_wdata_T_12 & _addr_aligned_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_dataMemory_out_en = io_in_mem_en & ~io_out_addr_misaligned; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 131:36]
  assign io_dataMemory_out_rlen = {{6'd0}, size}; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 132:27]
  assign io_dataMemory_out_wen = io_in_mem_en & io_in_info_op[3]; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 75:28]
  assign io_dataMemory_out_wstrb = req_wmask[7:0]; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 134:27]
  assign io_dataMemory_out_addr = io_in_mem_addr; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 135:27]
  assign io_dataMemory_out_wdata = _req_wdata_T_18 | _req_wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_addr_misaligned = io_in_mem_en & ~addr_aligned; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 140:35]
  assign io_out_access_fault = io_in_mem_en & io_dataMemory_in_access_fault; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 141:35]
  assign io_out_page_fault = io_in_mem_en & io_dataMemory_in_page_fault; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 142:35]
  assign io_out_rdata = partial_load ? rdata_partial_result : rdata64; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 139:32]
  assign io_out_ready = io_dataMemory_in_ready & io_dataMemory_out_en; // @[playground/src/pipeline/memory/lsu/LsExecute.scala 138:52]
endmodule
module Lsu(
  input         clock,
  input         reset,
  input         io_memoryUnit_in_mem_en, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [6:0]  io_memoryUnit_in_info_op, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_info_imm, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_info_inst, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_src_info_src1_data, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_src_info_src2_data, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_0, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_1, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_2, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_3, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_8, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_9, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_11, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_exception_12, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_0, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_1, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_2, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_3, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_4, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_5, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_6, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_7, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_8, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_9, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_10, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_ex_interrupt_11, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_ex_tval_0, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_ex_tval_1, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_ex_tval_2, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_ex_tval_12, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_lr, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_memoryUnit_in_lr_addr, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_memoryUnit_in_allow_to_go, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ready, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_rdata, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_0, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_1, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_2, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_3, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_4, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_5, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_6, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_7, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_8, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_9, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_11, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_12, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_13, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_exception_15, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_0, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_1, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_2, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_3, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_4, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_5, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_6, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_7, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_8, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_9, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_10, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_ex_interrupt_11, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_0, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_1, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_2, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_4, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_5, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_6, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_7, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_12, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_13, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_ex_tval_15, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_complete_single_request, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_lr_wen, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_memoryUnit_out_lr_wbit, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_memoryUnit_out_lr_waddr, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_dataMemory_in_access_fault, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_dataMemory_in_page_fault, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input         io_dataMemory_in_ready, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  input  [63:0] io_dataMemory_in_rdata, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_dataMemory_out_en, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [7:0]  io_dataMemory_out_rlen, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output        io_dataMemory_out_wen, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [7:0]  io_dataMemory_out_wstrb, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_dataMemory_out_addr, // @[playground/src/pipeline/memory/Lsu.scala 53:14]
  output [63:0] io_dataMemory_out_wdata // @[playground/src/pipeline/memory/Lsu.scala 53:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] AtomAlu_io_in_rdata; // @[playground/src/pipeline/memory/Lsu.scala 58:25]
  wire [63:0] AtomAlu_io_in_src2; // @[playground/src/pipeline/memory/Lsu.scala 58:25]
  wire [6:0] AtomAlu_io_in_info_op; // @[playground/src/pipeline/memory/Lsu.scala 58:25]
  wire [63:0] AtomAlu_io_in_info_inst; // @[playground/src/pipeline/memory/Lsu.scala 58:25]
  wire [63:0] AtomAlu_io_out_result; // @[playground/src/pipeline/memory/Lsu.scala 58:25]
  wire  LsExecute_io_dataMemory_in_access_fault; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_dataMemory_in_page_fault; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_dataMemory_in_ready; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [63:0] LsExecute_io_dataMemory_in_rdata; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_dataMemory_out_en; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [7:0] LsExecute_io_dataMemory_out_rlen; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_dataMemory_out_wen; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [7:0] LsExecute_io_dataMemory_out_wstrb; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [63:0] LsExecute_io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [63:0] LsExecute_io_dataMemory_out_wdata; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_in_mem_en; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [63:0] LsExecute_io_in_mem_addr; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [63:0] LsExecute_io_in_wdata; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [6:0] LsExecute_io_in_info_op; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_out_addr_misaligned; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_out_access_fault; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_out_page_fault; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire [63:0] LsExecute_io_out_rdata; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  LsExecute_io_out_ready; // @[playground/src/pipeline/memory/Lsu.scala 59:25]
  wire  store_req = io_memoryUnit_in_mem_en & io_memoryUnit_in_info_op[3]; // @[playground/src/pipeline/memory/Lsu.scala 68:25]
  wire  _load_req_T_4 = ~io_memoryUnit_in_info_op[3] & ~io_memoryUnit_in_info_op[5]; // @[playground/src/defines/isa/Instructions.scala 110:50]
  wire  load_req = io_memoryUnit_in_mem_en & _load_req_T_4; // @[playground/src/pipeline/memory/Lsu.scala 69:25]
  wire  atom_req = io_memoryUnit_in_mem_en & io_memoryUnit_in_info_op[5]; // @[playground/src/pipeline/memory/Lsu.scala 70:25]
  wire  _amo_req_T_1 = io_memoryUnit_in_info_op == 7'h20; // @[playground/src/defines/isa/Instructions.scala 111:40]
  wire  _amo_req_T_4 = io_memoryUnit_in_info_op == 7'h21; // @[playground/src/defines/isa/Instructions.scala 112:40]
  wire  _amo_req_T_6 = io_memoryUnit_in_info_op[5] & ~_amo_req_T_1 & ~_amo_req_T_4; // @[playground/src/defines/isa/Instructions.scala 113:63]
  wire  amo_req = io_memoryUnit_in_mem_en & _amo_req_T_6; // @[playground/src/pipeline/memory/Lsu.scala 71:25]
  wire  lr_req = io_memoryUnit_in_mem_en & _amo_req_T_1; // @[playground/src/pipeline/memory/Lsu.scala 72:25]
  wire  sc_req = io_memoryUnit_in_mem_en & _amo_req_T_4; // @[playground/src/pipeline/memory/Lsu.scala 73:25]
  wire [2:0] funct3 = io_memoryUnit_in_info_inst[14:12]; // @[playground/src/pipeline/memory/Lsu.scala 75:20]
  wire  atom_d = funct3[0]; // @[playground/src/pipeline/memory/Lsu.scala 76:22]
  reg [1:0] state; // @[playground/src/pipeline/memory/Lsu.scala 89:27]
  reg [63:0] atom_wdata; // @[playground/src/pipeline/memory/Lsu.scala 90:23]
  reg [63:0] atom_rdata; // @[playground/src/pipeline/memory/Lsu.scala 91:23]
  wire  sc_invalid = (io_memoryUnit_in_src_info_src1_data != io_memoryUnit_in_lr_addr | ~io_memoryUnit_in_lr) & sc_req; // @[playground/src/pipeline/memory/Lsu.scala 96:46]
  wire [63:0] _T_4 = io_memoryUnit_in_src_info_src1_data + io_memoryUnit_in_info_imm; // @[playground/src/pipeline/memory/Lsu.scala 114:39]
  wire [1:0] _T_5 = atom_d ? 2'h3 : 2'h2; // @[playground/src/pipeline/memory/Lsu.scala 121:39]
  wire [1:0] _GEN_0 = LsExecute_io_out_ready ? 2'h2 : state; // @[playground/src/pipeline/memory/Lsu.scala 124:35 125:17 89:27]
  wire  _GEN_1 = LsExecute_io_out_ready; // @[playground/src/pipeline/memory/Lsu.scala 107:27 124:35 127:35]
  wire  _GEN_2 = amo_req | io_memoryUnit_in_mem_en & ~atom_req; // @[playground/src/pipeline/memory/Lsu.scala 118:21 113:31 119:33]
  wire [63:0] _GEN_3 = amo_req ? io_memoryUnit_in_src_info_src1_data : _T_4; // @[playground/src/pipeline/memory/Lsu.scala 118:21 114:31 120:33]
  wire [6:0] _GEN_4 = amo_req ? {{5'd0}, _T_5} : io_memoryUnit_in_info_op; // @[playground/src/pipeline/memory/Lsu.scala 118:21 115:31 121:33]
  wire  _GEN_6 = amo_req ? 1'h0 : LsExecute_io_out_ready | sc_invalid; // @[playground/src/pipeline/memory/Lsu.scala 118:21 117:31 123:33]
  wire [1:0] _GEN_7 = amo_req ? _GEN_0 : state; // @[playground/src/pipeline/memory/Lsu.scala 118:21 89:27]
  wire  _GEN_8 = amo_req & _GEN_1; // @[playground/src/pipeline/memory/Lsu.scala 118:21 107:27]
  wire  _GEN_11 = lr_req | _GEN_2; // @[playground/src/pipeline/memory/Lsu.scala 132:20 133:33]
  wire [63:0] _GEN_12 = lr_req ? io_memoryUnit_in_src_info_src1_data : _GEN_3; // @[playground/src/pipeline/memory/Lsu.scala 132:20 134:33]
  wire [6:0] _GEN_13 = lr_req ? {{5'd0}, _T_5} : _GEN_4; // @[playground/src/pipeline/memory/Lsu.scala 132:20 135:33]
  wire  _GEN_15 = lr_req ? LsExecute_io_out_ready : _GEN_6; // @[playground/src/pipeline/memory/Lsu.scala 132:20 137:33]
  wire [1:0] _state_T = sc_invalid ? 2'h0 : 2'h1; // @[playground/src/pipeline/memory/Lsu.scala 139:34]
  wire [3:0] _T_8 = atom_d ? 4'hb : 4'ha; // @[playground/src/pipeline/memory/Lsu.scala 145:37]
  wire [1:0] _GEN_17 = io_memoryUnit_in_allow_to_go ? 2'h0 : state; // @[playground/src/pipeline/memory/Lsu.scala 148:25 149:15 89:27]
  wire  _GEN_22 = 2'h3 == state & LsExecute_io_out_ready; // @[playground/src/pipeline/memory/Lsu.scala 111:17 102:27 168:31]
  wire [1:0] _GEN_23 = 2'h3 == state ? _GEN_17 : state; // @[playground/src/pipeline/memory/Lsu.scala 111:17 89:27]
  wire  _GEN_24 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[playground/src/pipeline/memory/Lsu.scala 111:17 154:31]
  wire  _GEN_28 = 2'h2 == state ? 1'h0 : _GEN_22; // @[playground/src/pipeline/memory/Lsu.scala 111:17 158:31]
  wire [1:0] _GEN_29 = 2'h2 == state ? 2'h3 : _GEN_23; // @[playground/src/pipeline/memory/Lsu.scala 111:17 159:31]
  wire  _GEN_31 = 2'h1 == state | _GEN_24; // @[playground/src/pipeline/memory/Lsu.scala 111:17 143:31]
  wire [3:0] _GEN_33 = 2'h1 == state ? _T_8 : _T_8; // @[playground/src/pipeline/memory/Lsu.scala 111:17 145:31]
  wire [63:0] _GEN_34 = 2'h1 == state ? io_memoryUnit_in_src_info_src2_data : atom_wdata; // @[playground/src/pipeline/memory/Lsu.scala 111:17 146:31]
  wire  _GEN_35 = 2'h1 == state ? LsExecute_io_out_ready : _GEN_28; // @[playground/src/pipeline/memory/Lsu.scala 111:17 147:31]
  wire  _GEN_42 = 2'h0 == state ? _GEN_15 : _GEN_35; // @[playground/src/pipeline/memory/Lsu.scala 111:17]
  wire  _GEN_44 = 2'h0 == state & _GEN_8; // @[playground/src/pipeline/memory/Lsu.scala 111:17 107:27]
  wire  _T_12 = LsExecute_io_out_addr_misaligned | LsExecute_io_out_access_fault; // @[playground/src/pipeline/memory/Lsu.scala 176:35]
  wire  _T_13 = _T_12 | LsExecute_io_out_page_fault; // @[playground/src/pipeline/memory/Lsu.scala 177:34]
  wire  _io_memoryUnit_out_ex_exception_4_T = load_req | lr_req; // @[playground/src/pipeline/memory/Lsu.scala 188:67]
  wire  _io_memoryUnit_out_ex_exception_6_T_1 = store_req | sc_req | amo_req; // @[playground/src/pipeline/memory/Lsu.scala 192:76]
  wire [63:0] _io_memoryUnit_out_rdata_T = amo_req ? atom_rdata : LsExecute_io_out_rdata; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  AtomAlu AtomAlu ( // @[playground/src/pipeline/memory/Lsu.scala 58:25]
    .io_in_rdata(AtomAlu_io_in_rdata),
    .io_in_src2(AtomAlu_io_in_src2),
    .io_in_info_op(AtomAlu_io_in_info_op),
    .io_in_info_inst(AtomAlu_io_in_info_inst),
    .io_out_result(AtomAlu_io_out_result)
  );
  LsExecute LsExecute ( // @[playground/src/pipeline/memory/Lsu.scala 59:25]
    .io_dataMemory_in_access_fault(LsExecute_io_dataMemory_in_access_fault),
    .io_dataMemory_in_page_fault(LsExecute_io_dataMemory_in_page_fault),
    .io_dataMemory_in_ready(LsExecute_io_dataMemory_in_ready),
    .io_dataMemory_in_rdata(LsExecute_io_dataMemory_in_rdata),
    .io_dataMemory_out_en(LsExecute_io_dataMemory_out_en),
    .io_dataMemory_out_rlen(LsExecute_io_dataMemory_out_rlen),
    .io_dataMemory_out_wen(LsExecute_io_dataMemory_out_wen),
    .io_dataMemory_out_wstrb(LsExecute_io_dataMemory_out_wstrb),
    .io_dataMemory_out_addr(LsExecute_io_dataMemory_out_addr),
    .io_dataMemory_out_wdata(LsExecute_io_dataMemory_out_wdata),
    .io_in_mem_en(LsExecute_io_in_mem_en),
    .io_in_mem_addr(LsExecute_io_in_mem_addr),
    .io_in_wdata(LsExecute_io_in_wdata),
    .io_in_info_op(LsExecute_io_in_info_op),
    .io_out_addr_misaligned(LsExecute_io_out_addr_misaligned),
    .io_out_access_fault(LsExecute_io_out_access_fault),
    .io_out_page_fault(LsExecute_io_out_page_fault),
    .io_out_rdata(LsExecute_io_out_rdata),
    .io_out_ready(LsExecute_io_out_ready)
  );
  assign io_memoryUnit_out_ready = _T_13 | _GEN_42; // @[playground/src/pipeline/memory/Lsu.scala 179:5 181:29]
  assign io_memoryUnit_out_rdata = sc_req ? {{63'd0}, sc_invalid} : _io_memoryUnit_out_rdata_T; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  assign io_memoryUnit_out_ex_exception_0 = io_memoryUnit_in_ex_exception_0; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_1 = io_memoryUnit_in_ex_exception_1; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_2 = io_memoryUnit_in_ex_exception_2; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_3 = io_memoryUnit_in_ex_exception_3; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_4 = (load_req | lr_req) & LsExecute_io_out_addr_misaligned; // @[playground/src/pipeline/memory/Lsu.scala 188:78]
  assign io_memoryUnit_out_ex_exception_5 = _io_memoryUnit_out_ex_exception_4_T & LsExecute_io_out_access_fault; // @[playground/src/pipeline/memory/Lsu.scala 189:78]
  assign io_memoryUnit_out_ex_exception_6 = (store_req | sc_req | amo_req) & LsExecute_io_out_addr_misaligned; // @[playground/src/pipeline/memory/Lsu.scala 192:88]
  assign io_memoryUnit_out_ex_exception_7 = _io_memoryUnit_out_ex_exception_6_T_1 & LsExecute_io_out_addr_misaligned; // @[playground/src/pipeline/memory/Lsu.scala 193:88]
  assign io_memoryUnit_out_ex_exception_8 = io_memoryUnit_in_ex_exception_8; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_9 = io_memoryUnit_in_ex_exception_9; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_11 = io_memoryUnit_in_ex_exception_11; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_12 = io_memoryUnit_in_ex_exception_12; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_exception_13 = _io_memoryUnit_out_ex_exception_4_T & LsExecute_io_out_page_fault; // @[playground/src/pipeline/memory/Lsu.scala 190:78]
  assign io_memoryUnit_out_ex_exception_15 = _io_memoryUnit_out_ex_exception_6_T_1 & LsExecute_io_out_page_fault; // @[playground/src/pipeline/memory/Lsu.scala 194:88]
  assign io_memoryUnit_out_ex_interrupt_0 = io_memoryUnit_in_ex_interrupt_0; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_1 = io_memoryUnit_in_ex_interrupt_1; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_2 = io_memoryUnit_in_ex_interrupt_2; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_3 = io_memoryUnit_in_ex_interrupt_3; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_4 = io_memoryUnit_in_ex_interrupt_4; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_5 = io_memoryUnit_in_ex_interrupt_5; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_6 = io_memoryUnit_in_ex_interrupt_6; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_7 = io_memoryUnit_in_ex_interrupt_7; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_8 = io_memoryUnit_in_ex_interrupt_8; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_9 = io_memoryUnit_in_ex_interrupt_9; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_10 = io_memoryUnit_in_ex_interrupt_10; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_interrupt_11 = io_memoryUnit_in_ex_interrupt_11; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_tval_0 = io_memoryUnit_in_ex_tval_0; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_tval_1 = io_memoryUnit_in_ex_tval_1; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_tval_2 = io_memoryUnit_in_ex_tval_2; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_tval_4 = io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 196:50]
  assign io_memoryUnit_out_ex_tval_5 = io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 197:50]
  assign io_memoryUnit_out_ex_tval_6 = io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 199:50]
  assign io_memoryUnit_out_ex_tval_7 = io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 200:50]
  assign io_memoryUnit_out_ex_tval_12 = io_memoryUnit_in_ex_tval_12; // @[playground/src/pipeline/memory/Lsu.scala 187:54]
  assign io_memoryUnit_out_ex_tval_13 = io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 198:50]
  assign io_memoryUnit_out_ex_tval_15 = io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 201:50]
  assign io_memoryUnit_out_complete_single_request = _T_13 ? 1'h0 : _GEN_44; // @[playground/src/pipeline/memory/Lsu.scala 179:5 182:29]
  assign io_memoryUnit_out_lr_wen = io_memoryUnit_out_ready & (lr_req | sc_req); // @[playground/src/pipeline/memory/Lsu.scala 81:57]
  assign io_memoryUnit_out_lr_wbit = io_memoryUnit_in_mem_en & _amo_req_T_1; // @[playground/src/pipeline/memory/Lsu.scala 72:25]
  assign io_memoryUnit_out_lr_waddr = io_memoryUnit_in_src_info_src1_data; // @[playground/src/pipeline/memory/Lsu.scala 83:30]
  assign io_dataMemory_out_en = LsExecute_io_dataMemory_out_en; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign io_dataMemory_out_rlen = LsExecute_io_dataMemory_out_rlen; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign io_dataMemory_out_wen = LsExecute_io_dataMemory_out_wen; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign io_dataMemory_out_wstrb = LsExecute_io_dataMemory_out_wstrb; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign io_dataMemory_out_addr = LsExecute_io_dataMemory_out_addr; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign io_dataMemory_out_wdata = LsExecute_io_dataMemory_out_wdata; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign AtomAlu_io_in_rdata = atom_wdata; // @[playground/src/pipeline/memory/Lsu.scala 92:20]
  assign AtomAlu_io_in_src2 = io_memoryUnit_in_src_info_src2_data; // @[playground/src/pipeline/memory/Lsu.scala 93:20]
  assign AtomAlu_io_in_info_op = io_memoryUnit_in_info_op; // @[playground/src/pipeline/memory/Lsu.scala 94:20]
  assign AtomAlu_io_in_info_inst = io_memoryUnit_in_info_inst; // @[playground/src/pipeline/memory/Lsu.scala 94:20]
  assign LsExecute_io_dataMemory_in_access_fault = io_dataMemory_in_access_fault; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign LsExecute_io_dataMemory_in_page_fault = io_dataMemory_in_page_fault; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign LsExecute_io_dataMemory_in_ready = io_dataMemory_in_ready; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign LsExecute_io_dataMemory_in_rdata = io_dataMemory_in_rdata; // @[playground/src/pipeline/memory/Lsu.scala 185:17]
  assign LsExecute_io_in_mem_en = 2'h0 == state ? _GEN_11 : _GEN_31; // @[playground/src/pipeline/memory/Lsu.scala 111:17]
  assign LsExecute_io_in_mem_addr = 2'h0 == state ? _GEN_12 : io_memoryUnit_in_src_info_src1_data; // @[playground/src/pipeline/memory/Lsu.scala 111:17]
  assign LsExecute_io_in_wdata = 2'h0 == state ? io_memoryUnit_in_src_info_src2_data : _GEN_34; // @[playground/src/pipeline/memory/Lsu.scala 111:17]
  assign LsExecute_io_in_info_op = 2'h0 == state ? _GEN_13 : {{3'd0}, _GEN_33}; // @[playground/src/pipeline/memory/Lsu.scala 111:17]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/memory/Lsu.scala 89:27]
      state <= 2'h0; // @[playground/src/pipeline/memory/Lsu.scala 89:27]
    end else if (_T_13) begin // @[playground/src/pipeline/memory/Lsu.scala 179:5]
      state <= 2'h0; // @[playground/src/pipeline/memory/Lsu.scala 180:29]
    end else if (2'h0 == state) begin // @[playground/src/pipeline/memory/Lsu.scala 111:17]
      if (sc_req) begin // @[playground/src/pipeline/memory/Lsu.scala 139:20]
        state <= _state_T; // @[playground/src/pipeline/memory/Lsu.scala 139:28]
      end else begin
        state <= _GEN_7;
      end
    end else if (2'h1 == state) begin // @[playground/src/pipeline/memory/Lsu.scala 111:17]
      state <= _GEN_17;
    end else begin
      state <= _GEN_29;
    end
    if (2'h0 == state) begin // @[playground/src/pipeline/memory/Lsu.scala 111:17]
      if (amo_req) begin // @[playground/src/pipeline/memory/Lsu.scala 118:21]
        atom_wdata <= LsExecute_io_out_rdata; // @[playground/src/pipeline/memory/Lsu.scala 129:20]
      end
    end else if (!(2'h1 == state)) begin // @[playground/src/pipeline/memory/Lsu.scala 111:17]
      if (2'h2 == state) begin // @[playground/src/pipeline/memory/Lsu.scala 111:17]
        atom_wdata <= AtomAlu_io_out_result; // @[playground/src/pipeline/memory/Lsu.scala 160:31]
      end
    end
    if (2'h0 == state) begin // @[playground/src/pipeline/memory/Lsu.scala 111:17]
      if (amo_req) begin // @[playground/src/pipeline/memory/Lsu.scala 118:21]
        atom_rdata <= LsExecute_io_out_rdata; // @[playground/src/pipeline/memory/Lsu.scala 130:20]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  atom_wdata = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atom_rdata = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mou(
  input         io_in_info_valid, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  input  [2:0]  io_in_info_fusel, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  input  [6:0]  io_in_info_op, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  input  [63:0] io_in_pc, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  output        io_out_flush, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  output        io_out_fence_i, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  output        io_out_sfence_vma, // @[playground/src/pipeline/memory/Mou.scala 9:14]
  output [63:0] io_out_target // @[playground/src/pipeline/memory/Mou.scala 9:14]
);
  wire  valid = io_in_info_valid & io_in_info_fusel == 3'h4; // @[playground/src/pipeline/memory/Mou.scala 22:37]
  assign io_out_flush = io_in_info_valid & io_in_info_fusel == 3'h4; // @[playground/src/pipeline/memory/Mou.scala 22:37]
  assign io_out_fence_i = valid & io_in_info_op == 7'h1; // @[playground/src/pipeline/memory/Mou.scala 23:26]
  assign io_out_sfence_vma = valid & io_in_info_op == 7'h2; // @[playground/src/pipeline/memory/Mou.scala 24:26]
  assign io_out_target = io_in_pc + 64'h4; // @[playground/src/pipeline/memory/Mou.scala 29:33]
endmodule
module MemoryUnit(
  input         clock,
  input         reset,
  output        io_ctrl_flush, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_ctrl_mem_stall, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_ctrl_allow_to_go, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_ctrl_fence_i, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_ctrl_complete_single_request, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_ctrl_sfence_vma_valid, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_ctrl_sfence_vma_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_ctrl_sfence_vma_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_pc, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_info_valid, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [2:0]  io_memoryStage_inst_0_info_fusel, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [6:0]  io_memoryStage_inst_0_info_op, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_info_reg_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [4:0]  io_memoryStage_inst_0_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_info_imm, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_info_inst, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_exception_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_0_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_ex_tval_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_ex_tval_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_ex_tval_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_0_ex_tval_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_pc, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_info_valid, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [2:0]  io_memoryStage_inst_1_info_fusel, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [6:0]  io_memoryStage_inst_1_info_op, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_info_reg_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [4:0]  io_memoryStage_inst_1_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_info_imm, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_info_inst, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_src_info_src1_data, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_src_info_src2_data, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_exception_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_memoryStage_inst_1_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_ex_tval_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_ex_tval_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_ex_tval_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_memoryStage_inst_1_ex_tval_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_fetchUnit_flush, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_fetchUnit_target, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_decodeUnit_0_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [4:0]  io_decodeUnit_0_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_decodeUnit_0_wdata, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_decodeUnit_1_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [4:0]  io_decodeUnit_1_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_decodeUnit_1_wdata, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_pc, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_13, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_14, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_exception_15, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_13, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_14, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_ex_tval_15, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_info_valid, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [2:0]  io_csr_in_info_fusel, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [6:0]  io_csr_in_info_op, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_lr_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_csr_in_lr_wbit, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_csr_in_lr_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_csr_out_flush, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_csr_out_target, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_csr_out_lr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_csr_out_lr_addr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_pc, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_info_valid, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [2:0]  io_writeBackStage_inst_0_info_fusel, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_info_reg_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [4:0]  io_writeBackStage_inst_0_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_rd_info_wdata_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_rd_info_wdata_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_13, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_14, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_exception_15, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_0_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_13, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_14, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_0_ex_tval_15, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_pc, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_info_valid, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [2:0]  io_writeBackStage_inst_1_info_fusel, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_info_reg_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [4:0]  io_writeBackStage_inst_1_info_reg_waddr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_rd_info_wdata_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_rd_info_wdata_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_13, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_14, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_exception_15, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_writeBackStage_inst_1_ex_interrupt_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_0, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_1, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_2, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_3, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_4, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_5, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_6, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_7, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_8, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_9, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_10, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_11, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_12, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_13, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_14, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_writeBackStage_inst_1_ex_tval_15, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_dataMemory_in_access_fault, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_dataMemory_in_page_fault, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input         io_dataMemory_in_ready, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  input  [63:0] io_dataMemory_in_rdata, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_dataMemory_out_en, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [7:0]  io_dataMemory_out_rlen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output        io_dataMemory_out_wen, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [7:0]  io_dataMemory_out_wstrb, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_dataMemory_out_addr, // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
  output [63:0] io_dataMemory_out_wdata // @[playground/src/pipeline/memory/MemoryUnit.scala 13:14]
);
  wire  Lsu_clock; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_reset; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_mem_en; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [6:0] Lsu_io_memoryUnit_in_info_op; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_info_imm; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_info_inst; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_exception_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_ex_tval_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_ex_tval_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_ex_tval_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_ex_tval_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_lr; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_in_lr_addr; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_in_allow_to_go; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ready; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_rdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_13; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_exception_15; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_13; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_ex_tval_15; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_complete_single_request; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_lr_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_memoryUnit_out_lr_wbit; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_memoryUnit_out_lr_waddr; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_dataMemory_in_access_fault; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_dataMemory_in_page_fault; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_dataMemory_in_ready; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_dataMemory_in_rdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_dataMemory_out_en; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [7:0] Lsu_io_dataMemory_out_rlen; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Lsu_io_dataMemory_out_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [7:0] Lsu_io_dataMemory_out_wstrb; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_dataMemory_out_addr; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire [63:0] Lsu_io_dataMemory_out_wdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
  wire  Mou_io_in_info_valid; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire [2:0] Mou_io_in_info_fusel; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire [6:0] Mou_io_in_info_op; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire [63:0] Mou_io_in_pc; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire  Mou_io_out_flush; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire  Mou_io_out_fence_i; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire  Mou_io_out_sfence_vma; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire [63:0] Mou_io_out_target; // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
  wire  _lsu_sel_T = io_memoryStage_inst_0_info_fusel == 3'h1; // @[playground/src/pipeline/memory/MemoryUnit.scala 39:41]
  wire  _lsu_sel_T_1 = io_memoryStage_inst_0_info_valid & _lsu_sel_T; // @[playground/src/pipeline/memory/MemoryUnit.scala 38:39]
  wire [7:0] lsu_sel_lo = {4'h0,io_memoryStage_inst_0_ex_exception_3,io_memoryStage_inst_0_ex_exception_2,
    io_memoryStage_inst_0_ex_exception_1,io_memoryStage_inst_0_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _lsu_sel_T_2 = {2'h0,1'h0,io_memoryStage_inst_0_ex_exception_12,io_memoryStage_inst_0_ex_exception_11,1'h0
    ,io_memoryStage_inst_0_ex_exception_9,io_memoryStage_inst_0_ex_exception_8,lsu_sel_lo}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] lsu_sel_lo_1 = {io_memoryStage_inst_0_ex_interrupt_5,io_memoryStage_inst_0_ex_interrupt_4,
    io_memoryStage_inst_0_ex_interrupt_3,io_memoryStage_inst_0_ex_interrupt_2,io_memoryStage_inst_0_ex_interrupt_1,
    io_memoryStage_inst_0_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _lsu_sel_T_4 = {io_memoryStage_inst_0_ex_interrupt_11,io_memoryStage_inst_0_ex_interrupt_10,
    io_memoryStage_inst_0_ex_interrupt_9,io_memoryStage_inst_0_ex_interrupt_8,io_memoryStage_inst_0_ex_interrupt_7,
    io_memoryStage_inst_0_ex_interrupt_6,lsu_sel_lo_1}; // @[playground/src/defines/Util.scala 8:45]
  wire  _lsu_sel_T_6 = |_lsu_sel_T_2 | |_lsu_sel_T_4; // @[playground/src/defines/Util.scala 8:29]
  wire  _lsu_sel_T_7 = ~_lsu_sel_T_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 40:7]
  wire  lsu_sel_0 = _lsu_sel_T_1 & _lsu_sel_T_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 39:56]
  wire  _lsu_sel_T_9 = io_memoryStage_inst_1_info_fusel == 3'h1; // @[playground/src/pipeline/memory/MemoryUnit.scala 42:41]
  wire  _lsu_sel_T_10 = io_memoryStage_inst_1_info_valid & _lsu_sel_T_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 41:39]
  wire [7:0] lsu_sel_lo_2 = {4'h0,io_memoryStage_inst_1_ex_exception_3,io_memoryStage_inst_1_ex_exception_2,
    io_memoryStage_inst_1_ex_exception_1,io_memoryStage_inst_1_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _lsu_sel_T_11 = {2'h0,1'h0,io_memoryStage_inst_1_ex_exception_12,io_memoryStage_inst_1_ex_exception_11,1'h0
    ,io_memoryStage_inst_1_ex_exception_9,io_memoryStage_inst_1_ex_exception_8,lsu_sel_lo_2}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] lsu_sel_lo_3 = {io_memoryStage_inst_1_ex_interrupt_5,io_memoryStage_inst_1_ex_interrupt_4,
    io_memoryStage_inst_1_ex_interrupt_3,io_memoryStage_inst_1_ex_interrupt_2,io_memoryStage_inst_1_ex_interrupt_1,
    io_memoryStage_inst_1_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _lsu_sel_T_13 = {io_memoryStage_inst_1_ex_interrupt_11,io_memoryStage_inst_1_ex_interrupt_10,
    io_memoryStage_inst_1_ex_interrupt_9,io_memoryStage_inst_1_ex_interrupt_8,io_memoryStage_inst_1_ex_interrupt_7,
    io_memoryStage_inst_1_ex_interrupt_6,lsu_sel_lo_3}; // @[playground/src/defines/Util.scala 8:45]
  wire  _lsu_sel_T_15 = |_lsu_sel_T_11 | |_lsu_sel_T_13; // @[playground/src/defines/Util.scala 8:29]
  wire  _lsu_sel_T_16 = ~_lsu_sel_T_15; // @[playground/src/pipeline/memory/MemoryUnit.scala 43:7]
  wire  _lsu_sel_T_17 = _lsu_sel_T_10 & _lsu_sel_T_16; // @[playground/src/pipeline/memory/MemoryUnit.scala 42:56]
  wire  lsu_sel_1 = _lsu_sel_T_17 & _lsu_sel_T_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 43:45]
  wire [63:0] _T_1 = lsu_sel_0 ? io_memoryStage_inst_0_info_inst : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_2 = lsu_sel_1 ? io_memoryStage_inst_1_info_inst : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_4 = lsu_sel_0 ? io_memoryStage_inst_0_info_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_5 = lsu_sel_1 ? io_memoryStage_inst_1_info_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _T_13 = lsu_sel_0 ? io_memoryStage_inst_0_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _T_14 = lsu_sel_1 ? io_memoryStage_inst_1_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_37 = lsu_sel_0 ? io_memoryStage_inst_0_src_info_src2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_38 = lsu_sel_1 ? io_memoryStage_inst_1_src_info_src2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_40 = lsu_sel_0 ? io_memoryStage_inst_0_src_info_src1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_41 = lsu_sel_1 ? io_memoryStage_inst_1_src_info_src1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_43 = lsu_sel_0 ? io_memoryStage_inst_0_ex_tval_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_44 = lsu_sel_1 ? io_memoryStage_inst_1_ex_tval_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_46 = lsu_sel_0 ? io_memoryStage_inst_0_ex_tval_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_47 = lsu_sel_1 ? io_memoryStage_inst_1_ex_tval_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_49 = lsu_sel_0 ? io_memoryStage_inst_0_ex_tval_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_50 = lsu_sel_1 ? io_memoryStage_inst_1_ex_tval_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_79 = lsu_sel_0 ? io_memoryStage_inst_0_ex_tval_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _T_80 = lsu_sel_1 ? io_memoryStage_inst_1_ex_tval_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] csr_sel_lo = {io_writeBackStage_inst_0_ex_exception_7,io_writeBackStage_inst_0_ex_exception_6,
    io_writeBackStage_inst_0_ex_exception_5,io_writeBackStage_inst_0_ex_exception_4,
    io_writeBackStage_inst_0_ex_exception_3,io_writeBackStage_inst_0_ex_exception_2,
    io_writeBackStage_inst_0_ex_exception_1,io_writeBackStage_inst_0_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _csr_sel_T = {io_writeBackStage_inst_0_ex_exception_15,io_writeBackStage_inst_0_ex_exception_14,
    io_writeBackStage_inst_0_ex_exception_13,io_writeBackStage_inst_0_ex_exception_12,
    io_writeBackStage_inst_0_ex_exception_11,io_writeBackStage_inst_0_ex_exception_10,
    io_writeBackStage_inst_0_ex_exception_9,io_writeBackStage_inst_0_ex_exception_8,csr_sel_lo}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] csr_sel_lo_1 = {io_writeBackStage_inst_0_ex_interrupt_5,io_writeBackStage_inst_0_ex_interrupt_4,
    io_writeBackStage_inst_0_ex_interrupt_3,io_writeBackStage_inst_0_ex_interrupt_2,
    io_writeBackStage_inst_0_ex_interrupt_1,io_writeBackStage_inst_0_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _csr_sel_T_2 = {io_writeBackStage_inst_0_ex_interrupt_11,io_writeBackStage_inst_0_ex_interrupt_10,
    io_writeBackStage_inst_0_ex_interrupt_9,io_writeBackStage_inst_0_ex_interrupt_8,
    io_writeBackStage_inst_0_ex_interrupt_7,io_writeBackStage_inst_0_ex_interrupt_6,csr_sel_lo_1}; // @[playground/src/defines/Util.scala 8:45]
  wire  _csr_sel_T_4 = |_csr_sel_T | |_csr_sel_T_2; // @[playground/src/defines/Util.scala 8:29]
  wire [7:0] csr_sel_lo_2 = {io_writeBackStage_inst_1_ex_exception_7,io_writeBackStage_inst_1_ex_exception_6,
    io_writeBackStage_inst_1_ex_exception_5,io_writeBackStage_inst_1_ex_exception_4,
    io_writeBackStage_inst_1_ex_exception_3,io_writeBackStage_inst_1_ex_exception_2,
    io_writeBackStage_inst_1_ex_exception_1,io_writeBackStage_inst_1_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _csr_sel_T_5 = {io_writeBackStage_inst_1_ex_exception_15,io_writeBackStage_inst_1_ex_exception_14,
    io_writeBackStage_inst_1_ex_exception_13,io_writeBackStage_inst_1_ex_exception_12,
    io_writeBackStage_inst_1_ex_exception_11,io_writeBackStage_inst_1_ex_exception_10,
    io_writeBackStage_inst_1_ex_exception_9,io_writeBackStage_inst_1_ex_exception_8,csr_sel_lo_2}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] csr_sel_lo_3 = {io_writeBackStage_inst_1_ex_interrupt_5,io_writeBackStage_inst_1_ex_interrupt_4,
    io_writeBackStage_inst_1_ex_interrupt_3,io_writeBackStage_inst_1_ex_interrupt_2,
    io_writeBackStage_inst_1_ex_interrupt_1,io_writeBackStage_inst_1_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _csr_sel_T_7 = {io_writeBackStage_inst_1_ex_interrupt_11,io_writeBackStage_inst_1_ex_interrupt_10,
    io_writeBackStage_inst_1_ex_interrupt_9,io_writeBackStage_inst_1_ex_interrupt_8,
    io_writeBackStage_inst_1_ex_interrupt_7,io_writeBackStage_inst_1_ex_interrupt_6,csr_sel_lo_3}; // @[playground/src/defines/Util.scala 8:45]
  wire  _csr_sel_T_9 = |_csr_sel_T_5 | |_csr_sel_T_7; // @[playground/src/defines/Util.scala 8:29]
  wire  csr_sel = _csr_sel_T_4 | ~_csr_sel_T_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 53:45]
  wire  _io_csr_in_pc_T = ~csr_sel; // @[playground/src/pipeline/memory/MemoryUnit.scala 60:36]
  wire [63:0] _io_csr_in_pc_T_1 = csr_sel ? io_memoryStage_inst_0_pc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_pc_T_2 = _io_csr_in_pc_T ? io_memoryStage_inst_1_pc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_pc_T_3 = _io_csr_in_pc_T_1 | _io_csr_in_pc_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_1 = csr_sel ? io_writeBackStage_inst_0_ex_tval_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_2 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_3 = _io_csr_in_ex_T_1 | _io_csr_in_ex_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_4 = csr_sel ? io_writeBackStage_inst_0_ex_tval_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_5 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_6 = _io_csr_in_ex_T_4 | _io_csr_in_ex_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_7 = csr_sel ? io_writeBackStage_inst_0_ex_tval_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_8 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_9 = _io_csr_in_ex_T_7 | _io_csr_in_ex_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_10 = csr_sel ? io_writeBackStage_inst_0_ex_tval_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_11 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_12 = _io_csr_in_ex_T_10 | _io_csr_in_ex_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_13 = csr_sel ? io_writeBackStage_inst_0_ex_tval_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_14 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_15 = _io_csr_in_ex_T_13 | _io_csr_in_ex_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_16 = csr_sel ? io_writeBackStage_inst_0_ex_tval_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_17 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_18 = _io_csr_in_ex_T_16 | _io_csr_in_ex_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_19 = csr_sel ? io_writeBackStage_inst_0_ex_tval_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_20 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_21 = _io_csr_in_ex_T_19 | _io_csr_in_ex_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_22 = csr_sel ? io_writeBackStage_inst_0_ex_tval_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_23 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_24 = _io_csr_in_ex_T_22 | _io_csr_in_ex_T_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_25 = csr_sel ? io_writeBackStage_inst_0_ex_tval_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_26 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_27 = _io_csr_in_ex_T_25 | _io_csr_in_ex_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_28 = csr_sel ? io_writeBackStage_inst_0_ex_tval_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_29 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_30 = _io_csr_in_ex_T_28 | _io_csr_in_ex_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_31 = csr_sel ? io_writeBackStage_inst_0_ex_tval_10 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_32 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_10 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_33 = _io_csr_in_ex_T_31 | _io_csr_in_ex_T_32; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_34 = csr_sel ? io_writeBackStage_inst_0_ex_tval_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_35 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_36 = _io_csr_in_ex_T_34 | _io_csr_in_ex_T_35; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_37 = csr_sel ? io_writeBackStage_inst_0_ex_tval_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_38 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_39 = _io_csr_in_ex_T_37 | _io_csr_in_ex_T_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_40 = csr_sel ? io_writeBackStage_inst_0_ex_tval_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_41 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_42 = _io_csr_in_ex_T_40 | _io_csr_in_ex_T_41; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_43 = csr_sel ? io_writeBackStage_inst_0_ex_tval_14 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_44 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_14 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_45 = _io_csr_in_ex_T_43 | _io_csr_in_ex_T_44; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_46 = csr_sel ? io_writeBackStage_inst_0_ex_tval_15 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_47 = _io_csr_in_pc_T ? io_writeBackStage_inst_1_ex_tval_15 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_csr_in_ex_T_48 = _io_csr_in_ex_T_46 | _io_csr_in_ex_T_47; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_51 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_0 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_54 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_1 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_57 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_2 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_60 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_3 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_63 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_4 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_66 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_5 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_69 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_6 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_72 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_7 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_75 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_8 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_78 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_9 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_81 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_10 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_84 = csr_sel & io_writeBackStage_inst_0_ex_interrupt_11 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_interrupt_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_87 = csr_sel & io_writeBackStage_inst_0_ex_exception_0 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_90 = csr_sel & io_writeBackStage_inst_0_ex_exception_1 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_93 = csr_sel & io_writeBackStage_inst_0_ex_exception_2 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_96 = csr_sel & io_writeBackStage_inst_0_ex_exception_3 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_99 = csr_sel & io_writeBackStage_inst_0_ex_exception_4 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_102 = csr_sel & io_writeBackStage_inst_0_ex_exception_5 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_105 = csr_sel & io_writeBackStage_inst_0_ex_exception_6 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_108 = csr_sel & io_writeBackStage_inst_0_ex_exception_7 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_111 = csr_sel & io_writeBackStage_inst_0_ex_exception_8 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_114 = csr_sel & io_writeBackStage_inst_0_ex_exception_9 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_117 = csr_sel & io_writeBackStage_inst_0_ex_exception_10 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_120 = csr_sel & io_writeBackStage_inst_0_ex_exception_11 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_123 = csr_sel & io_writeBackStage_inst_0_ex_exception_12 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_126 = csr_sel & io_writeBackStage_inst_0_ex_exception_13 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_129 = csr_sel & io_writeBackStage_inst_0_ex_exception_14 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_ex_T_132 = csr_sel & io_writeBackStage_inst_0_ex_exception_15 | _io_csr_in_pc_T &
    io_writeBackStage_inst_1_ex_exception_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _io_csr_in_info_T_13 = csr_sel ? io_memoryStage_inst_0_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _io_csr_in_info_T_14 = _io_csr_in_pc_T ? io_memoryStage_inst_1_info_op : 7'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [6:0] _io_csr_in_info_T_15 = _io_csr_in_info_T_13 | _io_csr_in_info_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _io_csr_in_info_T_16 = csr_sel ? io_memoryStage_inst_0_info_fusel : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _io_csr_in_info_T_17 = _io_csr_in_pc_T ? io_memoryStage_inst_1_info_fusel : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _io_csr_in_info_T_18 = _io_csr_in_info_T_16 | _io_csr_in_info_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_csr_in_info_T_36 = csr_sel & io_memoryStage_inst_0_info_valid | _io_csr_in_pc_T &
    io_memoryStage_inst_1_info_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_58 = 3'h1 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_1 :
    io_writeBackStage_inst_0_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_59 = 3'h2 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_2 : _GEN_58
    ; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_60 = 3'h3 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_3 : _GEN_59
    ; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_61 = 3'h4 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_4 : _GEN_60
    ; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_64 = 3'h1 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_1 :
    io_writeBackStage_inst_1_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_65 = 3'h2 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_2 : _GEN_64
    ; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_66 = 3'h3 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_3 : _GEN_65
    ; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire [63:0] _GEN_67 = 3'h4 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_4 : _GEN_66
    ; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  wire  _io_writeBackStage_inst_1_info_valid_T_1 = ~(io_fetchUnit_flush & csr_sel); // @[playground/src/pipeline/memory/MemoryUnit.scala 92:5]
  Lsu Lsu ( // @[playground/src/pipeline/memory/MemoryUnit.scala 26:19]
    .clock(Lsu_clock),
    .reset(Lsu_reset),
    .io_memoryUnit_in_mem_en(Lsu_io_memoryUnit_in_mem_en),
    .io_memoryUnit_in_info_op(Lsu_io_memoryUnit_in_info_op),
    .io_memoryUnit_in_info_imm(Lsu_io_memoryUnit_in_info_imm),
    .io_memoryUnit_in_info_inst(Lsu_io_memoryUnit_in_info_inst),
    .io_memoryUnit_in_src_info_src1_data(Lsu_io_memoryUnit_in_src_info_src1_data),
    .io_memoryUnit_in_src_info_src2_data(Lsu_io_memoryUnit_in_src_info_src2_data),
    .io_memoryUnit_in_ex_exception_0(Lsu_io_memoryUnit_in_ex_exception_0),
    .io_memoryUnit_in_ex_exception_1(Lsu_io_memoryUnit_in_ex_exception_1),
    .io_memoryUnit_in_ex_exception_2(Lsu_io_memoryUnit_in_ex_exception_2),
    .io_memoryUnit_in_ex_exception_3(Lsu_io_memoryUnit_in_ex_exception_3),
    .io_memoryUnit_in_ex_exception_8(Lsu_io_memoryUnit_in_ex_exception_8),
    .io_memoryUnit_in_ex_exception_9(Lsu_io_memoryUnit_in_ex_exception_9),
    .io_memoryUnit_in_ex_exception_11(Lsu_io_memoryUnit_in_ex_exception_11),
    .io_memoryUnit_in_ex_exception_12(Lsu_io_memoryUnit_in_ex_exception_12),
    .io_memoryUnit_in_ex_interrupt_0(Lsu_io_memoryUnit_in_ex_interrupt_0),
    .io_memoryUnit_in_ex_interrupt_1(Lsu_io_memoryUnit_in_ex_interrupt_1),
    .io_memoryUnit_in_ex_interrupt_2(Lsu_io_memoryUnit_in_ex_interrupt_2),
    .io_memoryUnit_in_ex_interrupt_3(Lsu_io_memoryUnit_in_ex_interrupt_3),
    .io_memoryUnit_in_ex_interrupt_4(Lsu_io_memoryUnit_in_ex_interrupt_4),
    .io_memoryUnit_in_ex_interrupt_5(Lsu_io_memoryUnit_in_ex_interrupt_5),
    .io_memoryUnit_in_ex_interrupt_6(Lsu_io_memoryUnit_in_ex_interrupt_6),
    .io_memoryUnit_in_ex_interrupt_7(Lsu_io_memoryUnit_in_ex_interrupt_7),
    .io_memoryUnit_in_ex_interrupt_8(Lsu_io_memoryUnit_in_ex_interrupt_8),
    .io_memoryUnit_in_ex_interrupt_9(Lsu_io_memoryUnit_in_ex_interrupt_9),
    .io_memoryUnit_in_ex_interrupt_10(Lsu_io_memoryUnit_in_ex_interrupt_10),
    .io_memoryUnit_in_ex_interrupt_11(Lsu_io_memoryUnit_in_ex_interrupt_11),
    .io_memoryUnit_in_ex_tval_0(Lsu_io_memoryUnit_in_ex_tval_0),
    .io_memoryUnit_in_ex_tval_1(Lsu_io_memoryUnit_in_ex_tval_1),
    .io_memoryUnit_in_ex_tval_2(Lsu_io_memoryUnit_in_ex_tval_2),
    .io_memoryUnit_in_ex_tval_12(Lsu_io_memoryUnit_in_ex_tval_12),
    .io_memoryUnit_in_lr(Lsu_io_memoryUnit_in_lr),
    .io_memoryUnit_in_lr_addr(Lsu_io_memoryUnit_in_lr_addr),
    .io_memoryUnit_in_allow_to_go(Lsu_io_memoryUnit_in_allow_to_go),
    .io_memoryUnit_out_ready(Lsu_io_memoryUnit_out_ready),
    .io_memoryUnit_out_rdata(Lsu_io_memoryUnit_out_rdata),
    .io_memoryUnit_out_ex_exception_0(Lsu_io_memoryUnit_out_ex_exception_0),
    .io_memoryUnit_out_ex_exception_1(Lsu_io_memoryUnit_out_ex_exception_1),
    .io_memoryUnit_out_ex_exception_2(Lsu_io_memoryUnit_out_ex_exception_2),
    .io_memoryUnit_out_ex_exception_3(Lsu_io_memoryUnit_out_ex_exception_3),
    .io_memoryUnit_out_ex_exception_4(Lsu_io_memoryUnit_out_ex_exception_4),
    .io_memoryUnit_out_ex_exception_5(Lsu_io_memoryUnit_out_ex_exception_5),
    .io_memoryUnit_out_ex_exception_6(Lsu_io_memoryUnit_out_ex_exception_6),
    .io_memoryUnit_out_ex_exception_7(Lsu_io_memoryUnit_out_ex_exception_7),
    .io_memoryUnit_out_ex_exception_8(Lsu_io_memoryUnit_out_ex_exception_8),
    .io_memoryUnit_out_ex_exception_9(Lsu_io_memoryUnit_out_ex_exception_9),
    .io_memoryUnit_out_ex_exception_11(Lsu_io_memoryUnit_out_ex_exception_11),
    .io_memoryUnit_out_ex_exception_12(Lsu_io_memoryUnit_out_ex_exception_12),
    .io_memoryUnit_out_ex_exception_13(Lsu_io_memoryUnit_out_ex_exception_13),
    .io_memoryUnit_out_ex_exception_15(Lsu_io_memoryUnit_out_ex_exception_15),
    .io_memoryUnit_out_ex_interrupt_0(Lsu_io_memoryUnit_out_ex_interrupt_0),
    .io_memoryUnit_out_ex_interrupt_1(Lsu_io_memoryUnit_out_ex_interrupt_1),
    .io_memoryUnit_out_ex_interrupt_2(Lsu_io_memoryUnit_out_ex_interrupt_2),
    .io_memoryUnit_out_ex_interrupt_3(Lsu_io_memoryUnit_out_ex_interrupt_3),
    .io_memoryUnit_out_ex_interrupt_4(Lsu_io_memoryUnit_out_ex_interrupt_4),
    .io_memoryUnit_out_ex_interrupt_5(Lsu_io_memoryUnit_out_ex_interrupt_5),
    .io_memoryUnit_out_ex_interrupt_6(Lsu_io_memoryUnit_out_ex_interrupt_6),
    .io_memoryUnit_out_ex_interrupt_7(Lsu_io_memoryUnit_out_ex_interrupt_7),
    .io_memoryUnit_out_ex_interrupt_8(Lsu_io_memoryUnit_out_ex_interrupt_8),
    .io_memoryUnit_out_ex_interrupt_9(Lsu_io_memoryUnit_out_ex_interrupt_9),
    .io_memoryUnit_out_ex_interrupt_10(Lsu_io_memoryUnit_out_ex_interrupt_10),
    .io_memoryUnit_out_ex_interrupt_11(Lsu_io_memoryUnit_out_ex_interrupt_11),
    .io_memoryUnit_out_ex_tval_0(Lsu_io_memoryUnit_out_ex_tval_0),
    .io_memoryUnit_out_ex_tval_1(Lsu_io_memoryUnit_out_ex_tval_1),
    .io_memoryUnit_out_ex_tval_2(Lsu_io_memoryUnit_out_ex_tval_2),
    .io_memoryUnit_out_ex_tval_4(Lsu_io_memoryUnit_out_ex_tval_4),
    .io_memoryUnit_out_ex_tval_5(Lsu_io_memoryUnit_out_ex_tval_5),
    .io_memoryUnit_out_ex_tval_6(Lsu_io_memoryUnit_out_ex_tval_6),
    .io_memoryUnit_out_ex_tval_7(Lsu_io_memoryUnit_out_ex_tval_7),
    .io_memoryUnit_out_ex_tval_12(Lsu_io_memoryUnit_out_ex_tval_12),
    .io_memoryUnit_out_ex_tval_13(Lsu_io_memoryUnit_out_ex_tval_13),
    .io_memoryUnit_out_ex_tval_15(Lsu_io_memoryUnit_out_ex_tval_15),
    .io_memoryUnit_out_complete_single_request(Lsu_io_memoryUnit_out_complete_single_request),
    .io_memoryUnit_out_lr_wen(Lsu_io_memoryUnit_out_lr_wen),
    .io_memoryUnit_out_lr_wbit(Lsu_io_memoryUnit_out_lr_wbit),
    .io_memoryUnit_out_lr_waddr(Lsu_io_memoryUnit_out_lr_waddr),
    .io_dataMemory_in_access_fault(Lsu_io_dataMemory_in_access_fault),
    .io_dataMemory_in_page_fault(Lsu_io_dataMemory_in_page_fault),
    .io_dataMemory_in_ready(Lsu_io_dataMemory_in_ready),
    .io_dataMemory_in_rdata(Lsu_io_dataMemory_in_rdata),
    .io_dataMemory_out_en(Lsu_io_dataMemory_out_en),
    .io_dataMemory_out_rlen(Lsu_io_dataMemory_out_rlen),
    .io_dataMemory_out_wen(Lsu_io_dataMemory_out_wen),
    .io_dataMemory_out_wstrb(Lsu_io_dataMemory_out_wstrb),
    .io_dataMemory_out_addr(Lsu_io_dataMemory_out_addr),
    .io_dataMemory_out_wdata(Lsu_io_dataMemory_out_wdata)
  );
  Mou Mou ( // @[playground/src/pipeline/memory/MemoryUnit.scala 27:19]
    .io_in_info_valid(Mou_io_in_info_valid),
    .io_in_info_fusel(Mou_io_in_info_fusel),
    .io_in_info_op(Mou_io_in_info_op),
    .io_in_pc(Mou_io_in_pc),
    .io_out_flush(Mou_io_out_flush),
    .io_out_fence_i(Mou_io_out_fence_i),
    .io_out_sfence_vma(Mou_io_out_sfence_vma),
    .io_out_target(Mou_io_out_target)
  );
  assign io_ctrl_flush = io_fetchUnit_flush; // @[playground/src/pipeline/memory/MemoryUnit.scala 94:21]
  assign io_ctrl_mem_stall = ~Lsu_io_memoryUnit_out_ready & Lsu_io_memoryUnit_in_mem_en; // @[playground/src/pipeline/memory/MemoryUnit.scala 95:50]
  assign io_ctrl_fence_i = Mou_io_out_fence_i; // @[playground/src/pipeline/memory/MemoryUnit.scala 97:35]
  assign io_ctrl_complete_single_request = Lsu_io_memoryUnit_out_complete_single_request; // @[playground/src/pipeline/memory/MemoryUnit.scala 98:35]
  assign io_ctrl_sfence_vma_valid = Mou_io_out_sfence_vma; // @[playground/src/pipeline/memory/MemoryUnit.scala 100:31]
  assign io_ctrl_sfence_vma_src_info_src1_data = io_memoryStage_inst_0_src_info_src1_data; // @[playground/src/pipeline/memory/MemoryUnit.scala 101:31]
  assign io_ctrl_sfence_vma_src_info_src2_data = io_memoryStage_inst_0_src_info_src2_data; // @[playground/src/pipeline/memory/MemoryUnit.scala 101:31]
  assign io_fetchUnit_flush = io_ctrl_allow_to_go & (io_csr_out_flush | Mou_io_out_flush); // @[playground/src/pipeline/memory/MemoryUnit.scala 103:46]
  assign io_fetchUnit_target = io_csr_out_flush ? io_csr_out_target : Mou_io_out_target; // @[playground/src/pipeline/memory/MemoryUnit.scala 104:29]
  assign io_decodeUnit_0_wen = io_writeBackStage_inst_0_info_reg_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 76:28]
  assign io_decodeUnit_0_waddr = io_writeBackStage_inst_0_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryUnit.scala 77:28]
  assign io_decodeUnit_0_wdata = 3'h5 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_5
     : _GEN_61; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  assign io_decodeUnit_1_wen = io_writeBackStage_inst_1_info_reg_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 76:28]
  assign io_decodeUnit_1_waddr = io_writeBackStage_inst_1_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryUnit.scala 77:28]
  assign io_decodeUnit_1_wdata = 3'h5 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_5
     : _GEN_67; // @[playground/src/pipeline/memory/MemoryUnit.scala 78:{28,28}]
  assign io_csr_in_pc = io_ctrl_allow_to_go ? _io_csr_in_pc_T_3 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 55:18 63:29 64:20]
  assign io_csr_in_ex_exception_0 = io_ctrl_allow_to_go & _io_csr_in_ex_T_87; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_1 = io_ctrl_allow_to_go & _io_csr_in_ex_T_90; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_2 = io_ctrl_allow_to_go & _io_csr_in_ex_T_93; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_3 = io_ctrl_allow_to_go & _io_csr_in_ex_T_96; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_4 = io_ctrl_allow_to_go & _io_csr_in_ex_T_99; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_5 = io_ctrl_allow_to_go & _io_csr_in_ex_T_102; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_6 = io_ctrl_allow_to_go & _io_csr_in_ex_T_105; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_7 = io_ctrl_allow_to_go & _io_csr_in_ex_T_108; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_8 = io_ctrl_allow_to_go & _io_csr_in_ex_T_111; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_9 = io_ctrl_allow_to_go & _io_csr_in_ex_T_114; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_10 = io_ctrl_allow_to_go & _io_csr_in_ex_T_117; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_11 = io_ctrl_allow_to_go & _io_csr_in_ex_T_120; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_12 = io_ctrl_allow_to_go & _io_csr_in_ex_T_123; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_13 = io_ctrl_allow_to_go & _io_csr_in_ex_T_126; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_14 = io_ctrl_allow_to_go & _io_csr_in_ex_T_129; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_exception_15 = io_ctrl_allow_to_go & _io_csr_in_ex_T_132; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_0 = io_ctrl_allow_to_go & _io_csr_in_ex_T_51; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_1 = io_ctrl_allow_to_go & _io_csr_in_ex_T_54; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_2 = io_ctrl_allow_to_go & _io_csr_in_ex_T_57; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_3 = io_ctrl_allow_to_go & _io_csr_in_ex_T_60; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_4 = io_ctrl_allow_to_go & _io_csr_in_ex_T_63; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_5 = io_ctrl_allow_to_go & _io_csr_in_ex_T_66; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_6 = io_ctrl_allow_to_go & _io_csr_in_ex_T_69; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_7 = io_ctrl_allow_to_go & _io_csr_in_ex_T_72; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_8 = io_ctrl_allow_to_go & _io_csr_in_ex_T_75; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_9 = io_ctrl_allow_to_go & _io_csr_in_ex_T_78; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_10 = io_ctrl_allow_to_go & _io_csr_in_ex_T_81; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_interrupt_11 = io_ctrl_allow_to_go & _io_csr_in_ex_T_84; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_0 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_3 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_1 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_6 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_2 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_9 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_3 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_12 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_4 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_15 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_5 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_18 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_6 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_21 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_7 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_24 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_8 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_27 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_9 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_30 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_10 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_33 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_11 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_36 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_12 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_39 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_13 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_42 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_14 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_45 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_ex_tval_15 = io_ctrl_allow_to_go ? _io_csr_in_ex_T_48 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 56:18 63:29 65:20]
  assign io_csr_in_info_valid = io_ctrl_allow_to_go & _io_csr_in_info_T_36; // @[playground/src/pipeline/memory/MemoryUnit.scala 57:18 63:29 66:20]
  assign io_csr_in_info_fusel = io_ctrl_allow_to_go ? _io_csr_in_info_T_18 : 3'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 57:18 63:29 66:20]
  assign io_csr_in_info_op = io_ctrl_allow_to_go ? _io_csr_in_info_T_15 : 7'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 57:18 63:29 66:20]
  assign io_csr_in_lr_wen = Lsu_io_memoryUnit_out_lr_wen & io_ctrl_allow_to_go; // @[playground/src/pipeline/memory/MemoryUnit.scala 69:58]
  assign io_csr_in_lr_wbit = Lsu_io_memoryUnit_out_lr_wbit; // @[playground/src/pipeline/memory/MemoryUnit.scala 70:29]
  assign io_csr_in_lr_waddr = Lsu_io_memoryUnit_out_lr_waddr; // @[playground/src/pipeline/memory/MemoryUnit.scala 71:29]
  assign io_writeBackStage_inst_0_pc = io_memoryStage_inst_0_pc; // @[playground/src/pipeline/memory/MemoryUnit.scala 80:57]
  assign io_writeBackStage_inst_0_info_valid = io_memoryStage_inst_0_info_valid; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_0_info_fusel = io_memoryStage_inst_0_info_fusel; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_0_info_reg_wen = io_memoryStage_inst_0_info_reg_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_0_info_reg_waddr = io_memoryStage_inst_0_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_0_rd_info_wdata_0 = io_memoryStage_inst_0_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_0_rd_info_wdata_1 = Lsu_io_memoryUnit_out_rdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 83:57]
  assign io_writeBackStage_inst_0_rd_info_wdata_2 = io_memoryStage_inst_0_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_0_rd_info_wdata_3 = io_memoryStage_inst_0_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_0_rd_info_wdata_4 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_0_rd_info_wdata_5 = io_memoryStage_inst_0_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_0_ex_exception_0 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_0 :
    io_memoryStage_inst_0_ex_exception_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_1 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_1 :
    io_memoryStage_inst_0_ex_exception_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_2 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_2 :
    io_memoryStage_inst_0_ex_exception_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_3 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_3 :
    io_memoryStage_inst_0_ex_exception_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_4 = lsu_sel_0 & Lsu_io_memoryUnit_out_ex_exception_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_5 = lsu_sel_0 & Lsu_io_memoryUnit_out_ex_exception_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_6 = lsu_sel_0 & Lsu_io_memoryUnit_out_ex_exception_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_7 = lsu_sel_0 & Lsu_io_memoryUnit_out_ex_exception_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_8 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_8 :
    io_memoryStage_inst_0_ex_exception_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_9 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_9 :
    io_memoryStage_inst_0_ex_exception_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_10 = 1'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_11 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_11 :
    io_memoryStage_inst_0_ex_exception_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_12 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_exception_12 :
    io_memoryStage_inst_0_ex_exception_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_13 = lsu_sel_0 & Lsu_io_memoryUnit_out_ex_exception_13; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_14 = 1'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_exception_15 = lsu_sel_0 & Lsu_io_memoryUnit_out_ex_exception_15; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_0 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_0 :
    io_memoryStage_inst_0_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_1 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_1 :
    io_memoryStage_inst_0_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_2 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_2 :
    io_memoryStage_inst_0_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_3 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_3 :
    io_memoryStage_inst_0_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_4 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_4 :
    io_memoryStage_inst_0_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_5 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_5 :
    io_memoryStage_inst_0_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_6 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_6 :
    io_memoryStage_inst_0_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_7 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_7 :
    io_memoryStage_inst_0_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_8 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_8 :
    io_memoryStage_inst_0_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_9 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_9 :
    io_memoryStage_inst_0_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_10 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_10 :
    io_memoryStage_inst_0_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_interrupt_11 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_interrupt_11 :
    io_memoryStage_inst_0_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_0 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_0 :
    io_memoryStage_inst_0_ex_tval_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_1 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_1 :
    io_memoryStage_inst_0_ex_tval_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_2 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_2 :
    io_memoryStage_inst_0_ex_tval_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_3 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_4 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_4 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_5 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_5 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_6 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_6 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_7 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_7 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_8 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_9 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_10 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_11 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_12 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_12 :
    io_memoryStage_inst_0_ex_tval_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_13 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_13 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_14 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_0_ex_tval_15 = lsu_sel_0 ? Lsu_io_memoryUnit_out_ex_tval_15 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_pc = io_memoryStage_inst_1_pc; // @[playground/src/pipeline/memory/MemoryUnit.scala 80:57]
  assign io_writeBackStage_inst_1_info_valid = io_memoryStage_inst_1_info_valid &
    _io_writeBackStage_inst_1_info_valid_T_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 91:77]
  assign io_writeBackStage_inst_1_info_fusel = io_memoryStage_inst_1_info_fusel; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_1_info_reg_wen = io_memoryStage_inst_1_info_reg_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_1_info_reg_waddr = io_memoryStage_inst_1_info_reg_waddr; // @[playground/src/pipeline/memory/MemoryUnit.scala 81:57]
  assign io_writeBackStage_inst_1_rd_info_wdata_0 = io_memoryStage_inst_1_rd_info_wdata_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_1_rd_info_wdata_1 = Lsu_io_memoryUnit_out_rdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 83:57]
  assign io_writeBackStage_inst_1_rd_info_wdata_2 = io_memoryStage_inst_1_rd_info_wdata_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_1_rd_info_wdata_3 = io_memoryStage_inst_1_rd_info_wdata_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_1_rd_info_wdata_4 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_1_rd_info_wdata_5 = io_memoryStage_inst_1_rd_info_wdata_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 82:57]
  assign io_writeBackStage_inst_1_ex_exception_0 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_0 :
    io_memoryStage_inst_1_ex_exception_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_1 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_1 :
    io_memoryStage_inst_1_ex_exception_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_2 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_2 :
    io_memoryStage_inst_1_ex_exception_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_3 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_3 :
    io_memoryStage_inst_1_ex_exception_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_4 = lsu_sel_1 & Lsu_io_memoryUnit_out_ex_exception_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_5 = lsu_sel_1 & Lsu_io_memoryUnit_out_ex_exception_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_6 = lsu_sel_1 & Lsu_io_memoryUnit_out_ex_exception_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_7 = lsu_sel_1 & Lsu_io_memoryUnit_out_ex_exception_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_8 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_8 :
    io_memoryStage_inst_1_ex_exception_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_9 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_9 :
    io_memoryStage_inst_1_ex_exception_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_10 = 1'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_11 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_11 :
    io_memoryStage_inst_1_ex_exception_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_12 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_exception_12 :
    io_memoryStage_inst_1_ex_exception_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_13 = lsu_sel_1 & Lsu_io_memoryUnit_out_ex_exception_13; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_14 = 1'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_exception_15 = lsu_sel_1 & Lsu_io_memoryUnit_out_ex_exception_15; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_0 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_0 :
    io_memoryStage_inst_1_ex_interrupt_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_1 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_1 :
    io_memoryStage_inst_1_ex_interrupt_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_2 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_2 :
    io_memoryStage_inst_1_ex_interrupt_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_3 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_3 :
    io_memoryStage_inst_1_ex_interrupt_3; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_4 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_4 :
    io_memoryStage_inst_1_ex_interrupt_4; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_5 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_5 :
    io_memoryStage_inst_1_ex_interrupt_5; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_6 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_6 :
    io_memoryStage_inst_1_ex_interrupt_6; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_7 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_7 :
    io_memoryStage_inst_1_ex_interrupt_7; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_8 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_8 :
    io_memoryStage_inst_1_ex_interrupt_8; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_9 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_9 :
    io_memoryStage_inst_1_ex_interrupt_9; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_10 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_10 :
    io_memoryStage_inst_1_ex_interrupt_10; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_interrupt_11 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_interrupt_11 :
    io_memoryStage_inst_1_ex_interrupt_11; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_0 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_0 :
    io_memoryStage_inst_1_ex_tval_0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_1 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_1 :
    io_memoryStage_inst_1_ex_tval_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_2 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_2 :
    io_memoryStage_inst_1_ex_tval_2; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_3 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_4 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_4 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_5 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_5 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_6 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_6 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_7 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_7 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_8 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_9 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_10 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_11 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_12 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_12 :
    io_memoryStage_inst_1_ex_tval_12; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_13 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_13 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_14 = 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_writeBackStage_inst_1_ex_tval_15 = lsu_sel_1 ? Lsu_io_memoryUnit_out_ex_tval_15 : 64'h0; // @[playground/src/pipeline/memory/MemoryUnit.scala 84:40]
  assign io_dataMemory_out_en = Lsu_io_dataMemory_out_en; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign io_dataMemory_out_rlen = Lsu_io_dataMemory_out_rlen; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign io_dataMemory_out_wen = Lsu_io_dataMemory_out_wen; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign io_dataMemory_out_wstrb = Lsu_io_dataMemory_out_wstrb; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign io_dataMemory_out_addr = Lsu_io_dataMemory_out_addr; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign io_dataMemory_out_wdata = Lsu_io_dataMemory_out_wdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign Lsu_clock = clock;
  assign Lsu_reset = reset;
  assign Lsu_io_memoryUnit_in_mem_en = lsu_sel_0 | lsu_sel_1; // @[playground/src/pipeline/memory/MemoryUnit.scala 45:50]
  assign Lsu_io_memoryUnit_in_info_op = _T_13 | _T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_info_imm = _T_4 | _T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_info_inst = _T_1 | _T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_src_info_src1_data = _T_40 | _T_41; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_src_info_src2_data = _T_37 | _T_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_0 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_0 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_1 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_1 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_2 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_2 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_3 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_3 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_8 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_8 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_9 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_9 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_11 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_11 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_exception_12 = lsu_sel_0 & io_memoryStage_inst_0_ex_exception_12 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_exception_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_0 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_0 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_1 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_1 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_2 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_2 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_3 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_3 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_4 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_4 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_5 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_5 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_6 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_6 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_7 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_7 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_8 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_8 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_9 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_9 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_10 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_10 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_interrupt_11 = lsu_sel_0 & io_memoryStage_inst_0_ex_interrupt_11 | lsu_sel_1 &
    io_memoryStage_inst_1_ex_interrupt_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_tval_0 = _T_43 | _T_44; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_tval_1 = _T_46 | _T_47; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_tval_2 = _T_49 | _T_50; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_ex_tval_12 = _T_79 | _T_80; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign Lsu_io_memoryUnit_in_lr = io_csr_out_lr; // @[playground/src/pipeline/memory/MemoryUnit.scala 72:29]
  assign Lsu_io_memoryUnit_in_lr_addr = io_csr_out_lr_addr; // @[playground/src/pipeline/memory/MemoryUnit.scala 73:29]
  assign Lsu_io_memoryUnit_in_allow_to_go = io_ctrl_allow_to_go; // @[playground/src/pipeline/memory/MemoryUnit.scala 50:33]
  assign Lsu_io_dataMemory_in_access_fault = io_dataMemory_in_access_fault; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign Lsu_io_dataMemory_in_page_fault = io_dataMemory_in_page_fault; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign Lsu_io_dataMemory_in_ready = io_dataMemory_in_ready; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign Lsu_io_dataMemory_in_rdata = io_dataMemory_in_rdata; // @[playground/src/pipeline/memory/MemoryUnit.scala 49:18]
  assign Mou_io_in_info_valid = io_memoryStage_inst_0_info_valid; // @[playground/src/pipeline/memory/MemoryUnit.scala 29:15]
  assign Mou_io_in_info_fusel = io_memoryStage_inst_0_info_fusel; // @[playground/src/pipeline/memory/MemoryUnit.scala 29:15]
  assign Mou_io_in_info_op = io_memoryStage_inst_0_info_op; // @[playground/src/pipeline/memory/MemoryUnit.scala 29:15]
  assign Mou_io_in_pc = io_memoryStage_inst_0_pc; // @[playground/src/pipeline/memory/MemoryUnit.scala 30:15]
endmodule
module WriteBackStage(
  input         clock,
  input         reset,
  input         io_ctrl_allow_to_go, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_0_pc, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_info_valid, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [2:0]  io_memoryUnit_inst_0_info_fusel, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_info_reg_wen, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [4:0]  io_memoryUnit_inst_0_info_reg_waddr, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_0_rd_info_wdata_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_12, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_13, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_exception_15, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_10, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_0_ex_interrupt_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_1_pc, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_info_valid, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [2:0]  io_memoryUnit_inst_1_info_fusel, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_info_reg_wen, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [4:0]  io_memoryUnit_inst_1_info_reg_waddr, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_1_rd_info_wdata_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input  [63:0] io_memoryUnit_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_12, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_13, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_exception_15, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_10, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  input         io_memoryUnit_inst_1_ex_interrupt_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_0_pc, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_info_valid, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [2:0]  io_writeBackUnit_inst_0_info_fusel, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_info_reg_wen, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [4:0]  io_writeBackUnit_inst_0_info_reg_waddr, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_0_rd_info_wdata_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_12, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_13, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_exception_15, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_10, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_0_ex_interrupt_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_1_pc, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_info_valid, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [2:0]  io_writeBackUnit_inst_1_info_fusel, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_info_reg_wen, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [4:0]  io_writeBackUnit_inst_1_info_reg_waddr, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_1_rd_info_wdata_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output [63:0] io_writeBackUnit_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_11, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_12, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_13, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_exception_15, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_0, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_1, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_2, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_3, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_4, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_5, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_6, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_7, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_8, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_9, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_10, // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
  output        io_writeBackUnit_inst_1_ex_interrupt_11 // @[playground/src/pipeline/writeback/WriteBackStage.scala 20:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] inst_0_pc; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_info_valid; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [2:0] inst_0_info_fusel; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [4:0] inst_0_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_0_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_0_rd_info_wdata_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_0_rd_info_wdata_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_0_rd_info_wdata_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_0_rd_info_wdata_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_12; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_13; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_exception_15; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_10; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_0_ex_interrupt_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_1_pc; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_info_valid; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [2:0] inst_1_info_fusel; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [4:0] inst_1_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_1_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_1_rd_info_wdata_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_1_rd_info_wdata_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_1_rd_info_wdata_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg [63:0] inst_1_rd_info_wdata_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_12; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_13; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_exception_15; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_10; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  reg  inst_1_ex_interrupt_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
  assign io_writeBackUnit_inst_0_pc = inst_0_pc; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_info_valid = inst_0_info_valid; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_info_fusel = inst_0_info_fusel; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_info_reg_wen = inst_0_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_info_reg_waddr = inst_0_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_rd_info_wdata_0 = inst_0_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_rd_info_wdata_1 = inst_0_rd_info_wdata_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_rd_info_wdata_2 = inst_0_rd_info_wdata_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_rd_info_wdata_3 = inst_0_rd_info_wdata_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_rd_info_wdata_5 = inst_0_rd_info_wdata_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_0 = inst_0_ex_exception_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_1 = inst_0_ex_exception_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_2 = inst_0_ex_exception_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_3 = inst_0_ex_exception_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_4 = inst_0_ex_exception_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_5 = inst_0_ex_exception_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_6 = inst_0_ex_exception_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_7 = inst_0_ex_exception_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_8 = inst_0_ex_exception_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_9 = inst_0_ex_exception_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_11 = inst_0_ex_exception_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_12 = inst_0_ex_exception_12; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_13 = inst_0_ex_exception_13; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_exception_15 = inst_0_ex_exception_15; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_0 = inst_0_ex_interrupt_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_1 = inst_0_ex_interrupt_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_2 = inst_0_ex_interrupt_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_3 = inst_0_ex_interrupt_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_4 = inst_0_ex_interrupt_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_5 = inst_0_ex_interrupt_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_6 = inst_0_ex_interrupt_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_7 = inst_0_ex_interrupt_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_8 = inst_0_ex_interrupt_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_9 = inst_0_ex_interrupt_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_10 = inst_0_ex_interrupt_10; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_0_ex_interrupt_11 = inst_0_ex_interrupt_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_pc = inst_1_pc; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_info_valid = inst_1_info_valid; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_info_fusel = inst_1_info_fusel; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_info_reg_wen = inst_1_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_info_reg_waddr = inst_1_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_rd_info_wdata_0 = inst_1_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_rd_info_wdata_1 = inst_1_rd_info_wdata_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_rd_info_wdata_2 = inst_1_rd_info_wdata_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_rd_info_wdata_3 = inst_1_rd_info_wdata_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_rd_info_wdata_5 = inst_1_rd_info_wdata_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_0 = inst_1_ex_exception_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_1 = inst_1_ex_exception_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_2 = inst_1_ex_exception_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_3 = inst_1_ex_exception_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_4 = inst_1_ex_exception_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_5 = inst_1_ex_exception_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_6 = inst_1_ex_exception_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_7 = inst_1_ex_exception_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_8 = inst_1_ex_exception_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_9 = inst_1_ex_exception_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_11 = inst_1_ex_exception_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_12 = inst_1_ex_exception_12; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_13 = inst_1_ex_exception_13; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_exception_15 = inst_1_ex_exception_15; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_0 = inst_1_ex_interrupt_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_1 = inst_1_ex_interrupt_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_2 = inst_1_ex_interrupt_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_3 = inst_1_ex_interrupt_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_4 = inst_1_ex_interrupt_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_5 = inst_1_ex_interrupt_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_6 = inst_1_ex_interrupt_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_7 = inst_1_ex_interrupt_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_8 = inst_1_ex_interrupt_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_9 = inst_1_ex_interrupt_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_10 = inst_1_ex_interrupt_10; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  assign io_writeBackUnit_inst_1_ex_interrupt_11 = inst_1_ex_interrupt_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 39:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_pc <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_pc <= io_memoryUnit_inst_0_pc; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_info_valid <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_info_valid <= io_memoryUnit_inst_0_info_valid; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_info_fusel <= 3'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_info_fusel <= io_memoryUnit_inst_0_info_fusel; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_info_reg_wen <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_info_reg_wen <= io_memoryUnit_inst_0_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_info_reg_waddr <= io_memoryUnit_inst_0_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_rd_info_wdata_0 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_rd_info_wdata_0 <= io_memoryUnit_inst_0_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_rd_info_wdata_1 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_rd_info_wdata_1 <= io_memoryUnit_inst_0_rd_info_wdata_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_rd_info_wdata_2 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_rd_info_wdata_2 <= io_memoryUnit_inst_0_rd_info_wdata_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_rd_info_wdata_3 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_rd_info_wdata_3 <= io_memoryUnit_inst_0_rd_info_wdata_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_rd_info_wdata_5 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_rd_info_wdata_5 <= io_memoryUnit_inst_0_rd_info_wdata_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_0 <= io_memoryUnit_inst_0_ex_exception_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_1 <= io_memoryUnit_inst_0_ex_exception_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_2 <= io_memoryUnit_inst_0_ex_exception_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_3 <= io_memoryUnit_inst_0_ex_exception_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_4 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_4 <= io_memoryUnit_inst_0_ex_exception_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_5 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_5 <= io_memoryUnit_inst_0_ex_exception_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_6 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_6 <= io_memoryUnit_inst_0_ex_exception_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_7 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_7 <= io_memoryUnit_inst_0_ex_exception_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_8 <= io_memoryUnit_inst_0_ex_exception_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_9 <= io_memoryUnit_inst_0_ex_exception_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_11 <= io_memoryUnit_inst_0_ex_exception_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_12 <= io_memoryUnit_inst_0_ex_exception_12; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_13 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_13 <= io_memoryUnit_inst_0_ex_exception_13; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_exception_15 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_exception_15 <= io_memoryUnit_inst_0_ex_exception_15; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_0 <= io_memoryUnit_inst_0_ex_interrupt_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_1 <= io_memoryUnit_inst_0_ex_interrupt_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_2 <= io_memoryUnit_inst_0_ex_interrupt_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_3 <= io_memoryUnit_inst_0_ex_interrupt_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_4 <= io_memoryUnit_inst_0_ex_interrupt_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_5 <= io_memoryUnit_inst_0_ex_interrupt_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_6 <= io_memoryUnit_inst_0_ex_interrupt_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_7 <= io_memoryUnit_inst_0_ex_interrupt_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_8 <= io_memoryUnit_inst_0_ex_interrupt_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_9 <= io_memoryUnit_inst_0_ex_interrupt_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_10 <= io_memoryUnit_inst_0_ex_interrupt_10; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_0_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_0_ex_interrupt_11 <= io_memoryUnit_inst_0_ex_interrupt_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_pc <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_pc <= io_memoryUnit_inst_1_pc; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_info_valid <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_info_valid <= io_memoryUnit_inst_1_info_valid; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_info_fusel <= 3'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_info_fusel <= io_memoryUnit_inst_1_info_fusel; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_info_reg_wen <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_info_reg_wen <= io_memoryUnit_inst_1_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_info_reg_waddr <= 5'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_info_reg_waddr <= io_memoryUnit_inst_1_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_rd_info_wdata_0 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_rd_info_wdata_0 <= io_memoryUnit_inst_1_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_rd_info_wdata_1 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_rd_info_wdata_1 <= io_memoryUnit_inst_1_rd_info_wdata_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_rd_info_wdata_2 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_rd_info_wdata_2 <= io_memoryUnit_inst_1_rd_info_wdata_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_rd_info_wdata_3 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_rd_info_wdata_3 <= io_memoryUnit_inst_1_rd_info_wdata_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_rd_info_wdata_5 <= 64'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_rd_info_wdata_5 <= io_memoryUnit_inst_1_rd_info_wdata_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_0 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_0 <= io_memoryUnit_inst_1_ex_exception_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_1 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_1 <= io_memoryUnit_inst_1_ex_exception_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_2 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_2 <= io_memoryUnit_inst_1_ex_exception_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_3 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_3 <= io_memoryUnit_inst_1_ex_exception_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_4 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_4 <= io_memoryUnit_inst_1_ex_exception_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_5 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_5 <= io_memoryUnit_inst_1_ex_exception_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_6 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_6 <= io_memoryUnit_inst_1_ex_exception_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_7 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_7 <= io_memoryUnit_inst_1_ex_exception_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_8 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_8 <= io_memoryUnit_inst_1_ex_exception_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_9 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_9 <= io_memoryUnit_inst_1_ex_exception_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_11 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_11 <= io_memoryUnit_inst_1_ex_exception_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_12 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_12 <= io_memoryUnit_inst_1_ex_exception_12; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_13 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_13 <= io_memoryUnit_inst_1_ex_exception_13; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_exception_15 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_exception_15 <= io_memoryUnit_inst_1_ex_exception_15; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_0 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_0 <= io_memoryUnit_inst_1_ex_interrupt_0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_1 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_1 <= io_memoryUnit_inst_1_ex_interrupt_1; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_2 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_2 <= io_memoryUnit_inst_1_ex_interrupt_2; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_3 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_3 <= io_memoryUnit_inst_1_ex_interrupt_3; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_4 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_4 <= io_memoryUnit_inst_1_ex_interrupt_4; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_5 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_5 <= io_memoryUnit_inst_1_ex_interrupt_5; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_6 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_6 <= io_memoryUnit_inst_1_ex_interrupt_6; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_7 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_7 <= io_memoryUnit_inst_1_ex_interrupt_7; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_8 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_8 <= io_memoryUnit_inst_1_ex_interrupt_8; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_9 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_9 <= io_memoryUnit_inst_1_ex_interrupt_9; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_10 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_10 <= io_memoryUnit_inst_1_ex_interrupt_10; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
    if (reset) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
      inst_1_ex_interrupt_11 <= 1'h0; // @[playground/src/pipeline/writeback/WriteBackStage.scala 29:51]
    end else if (io_ctrl_allow_to_go) begin // @[playground/src/pipeline/writeback/WriteBackStage.scala 34:37]
      inst_1_ex_interrupt_11 <= io_memoryUnit_inst_1_ex_interrupt_11; // @[playground/src/pipeline/writeback/WriteBackStage.scala 35:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  inst_0_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  inst_0_info_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_0_info_fusel = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  inst_0_info_reg_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  inst_0_info_reg_waddr = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  inst_0_rd_info_wdata_0 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  inst_0_rd_info_wdata_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  inst_0_rd_info_wdata_2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  inst_0_rd_info_wdata_3 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  inst_0_rd_info_wdata_5 = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  inst_0_ex_exception_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inst_0_ex_exception_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inst_0_ex_exception_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inst_0_ex_exception_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inst_0_ex_exception_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inst_0_ex_exception_5 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  inst_0_ex_exception_6 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  inst_0_ex_exception_7 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  inst_0_ex_exception_8 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  inst_0_ex_exception_9 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inst_0_ex_exception_11 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  inst_0_ex_exception_12 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  inst_0_ex_exception_13 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  inst_0_ex_exception_15 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  inst_0_ex_interrupt_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  inst_0_ex_interrupt_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  inst_0_ex_interrupt_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  inst_0_ex_interrupt_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  inst_0_ex_interrupt_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inst_0_ex_interrupt_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  inst_0_ex_interrupt_6 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  inst_0_ex_interrupt_7 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  inst_0_ex_interrupt_8 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  inst_0_ex_interrupt_9 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  inst_0_ex_interrupt_10 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  inst_0_ex_interrupt_11 = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  inst_1_pc = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  inst_1_info_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  inst_1_info_fusel = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  inst_1_info_reg_wen = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  inst_1_info_reg_waddr = _RAND_40[4:0];
  _RAND_41 = {2{`RANDOM}};
  inst_1_rd_info_wdata_0 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  inst_1_rd_info_wdata_1 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  inst_1_rd_info_wdata_2 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  inst_1_rd_info_wdata_3 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  inst_1_rd_info_wdata_5 = _RAND_45[63:0];
  _RAND_46 = {1{`RANDOM}};
  inst_1_ex_exception_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  inst_1_ex_exception_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  inst_1_ex_exception_2 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  inst_1_ex_exception_3 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  inst_1_ex_exception_4 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  inst_1_ex_exception_5 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  inst_1_ex_exception_6 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  inst_1_ex_exception_7 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  inst_1_ex_exception_8 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  inst_1_ex_exception_9 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  inst_1_ex_exception_11 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  inst_1_ex_exception_12 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  inst_1_ex_exception_13 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  inst_1_ex_exception_15 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  inst_1_ex_interrupt_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  inst_1_ex_interrupt_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  inst_1_ex_interrupt_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  inst_1_ex_interrupt_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  inst_1_ex_interrupt_4 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  inst_1_ex_interrupt_5 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  inst_1_ex_interrupt_6 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  inst_1_ex_interrupt_7 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  inst_1_ex_interrupt_8 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  inst_1_ex_interrupt_9 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  inst_1_ex_interrupt_10 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  inst_1_ex_interrupt_11 = _RAND_71[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBackUnit(
  input         clock,
  input         io_ctrl_allow_to_go, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_0_pc, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_info_valid, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [2:0]  io_writeBackStage_inst_0_info_fusel, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_info_reg_wen, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [4:0]  io_writeBackStage_inst_0_info_reg_waddr, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_0_rd_info_wdata_0, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_0_rd_info_wdata_1, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_0_rd_info_wdata_2, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_0_rd_info_wdata_3, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_0_rd_info_wdata_5, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_0, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_1, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_2, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_3, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_4, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_5, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_6, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_7, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_8, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_9, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_11, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_12, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_13, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_exception_15, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_0, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_1, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_2, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_3, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_4, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_5, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_6, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_7, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_8, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_9, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_10, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_0_ex_interrupt_11, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_1_pc, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_info_valid, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [2:0]  io_writeBackStage_inst_1_info_fusel, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_info_reg_wen, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [4:0]  io_writeBackStage_inst_1_info_reg_waddr, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_1_rd_info_wdata_0, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_1_rd_info_wdata_1, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_1_rd_info_wdata_2, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_1_rd_info_wdata_3, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input  [63:0] io_writeBackStage_inst_1_rd_info_wdata_5, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_0, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_1, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_2, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_3, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_4, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_5, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_6, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_7, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_8, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_9, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_11, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_12, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_13, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_exception_15, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_0, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_1, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_2, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_3, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_4, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_5, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_6, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_7, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_8, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_9, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_10, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  input         io_writeBackStage_inst_1_ex_interrupt_11, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output        io_regfile_0_wen, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [4:0]  io_regfile_0_waddr, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [63:0] io_regfile_0_wdata, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output        io_regfile_1_wen, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [4:0]  io_regfile_1_waddr, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [63:0] io_regfile_1_wdata, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [63:0] io_debug_wb_pc, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output        io_debug_wb_rf_wen, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [4:0]  io_debug_wb_rf_wnum, // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
  output [63:0] io_debug_wb_rf_wdata // @[playground/src/pipeline/writeback/WriteBackUnit.scala 11:14]
);
  wire  _io_regfile_0_wen_T = io_writeBackStage_inst_0_info_valid & io_writeBackStage_inst_0_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 19:42]
  wire  _io_regfile_0_wen_T_1 = _io_regfile_0_wen_T & io_ctrl_allow_to_go; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 20:46]
  wire [7:0] io_regfile_0_wen_lo = {io_writeBackStage_inst_0_ex_exception_7,io_writeBackStage_inst_0_ex_exception_6,
    io_writeBackStage_inst_0_ex_exception_5,io_writeBackStage_inst_0_ex_exception_4,
    io_writeBackStage_inst_0_ex_exception_3,io_writeBackStage_inst_0_ex_exception_2,
    io_writeBackStage_inst_0_ex_exception_1,io_writeBackStage_inst_0_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _io_regfile_0_wen_T_2 = {io_writeBackStage_inst_0_ex_exception_15,1'h0,
    io_writeBackStage_inst_0_ex_exception_13,io_writeBackStage_inst_0_ex_exception_12,
    io_writeBackStage_inst_0_ex_exception_11,1'h0,io_writeBackStage_inst_0_ex_exception_9,
    io_writeBackStage_inst_0_ex_exception_8,io_regfile_0_wen_lo}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] io_regfile_0_wen_lo_1 = {io_writeBackStage_inst_0_ex_interrupt_5,io_writeBackStage_inst_0_ex_interrupt_4,
    io_writeBackStage_inst_0_ex_interrupt_3,io_writeBackStage_inst_0_ex_interrupt_2,
    io_writeBackStage_inst_0_ex_interrupt_1,io_writeBackStage_inst_0_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _io_regfile_0_wen_T_4 = {io_writeBackStage_inst_0_ex_interrupt_11,io_writeBackStage_inst_0_ex_interrupt_10
    ,io_writeBackStage_inst_0_ex_interrupt_9,io_writeBackStage_inst_0_ex_interrupt_8,
    io_writeBackStage_inst_0_ex_interrupt_7,io_writeBackStage_inst_0_ex_interrupt_6,io_regfile_0_wen_lo_1}; // @[playground/src/defines/Util.scala 8:45]
  wire  _io_regfile_0_wen_T_6 = |_io_regfile_0_wen_T_2 | |_io_regfile_0_wen_T_4; // @[playground/src/defines/Util.scala 8:29]
  wire  _io_regfile_0_wen_T_7 = ~_io_regfile_0_wen_T_6; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 22:7]
  wire  _io_regfile_1_wen_T = io_writeBackStage_inst_1_info_valid & io_writeBackStage_inst_1_info_reg_wen; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 25:42]
  wire  _io_regfile_1_wen_T_1 = _io_regfile_1_wen_T & io_ctrl_allow_to_go; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 26:46]
  wire  _io_regfile_1_wen_T_8 = _io_regfile_1_wen_T_1 & _io_regfile_0_wen_T_7; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 27:27]
  wire [7:0] io_regfile_1_wen_lo_2 = {io_writeBackStage_inst_1_ex_exception_7,io_writeBackStage_inst_1_ex_exception_6,
    io_writeBackStage_inst_1_ex_exception_5,io_writeBackStage_inst_1_ex_exception_4,
    io_writeBackStage_inst_1_ex_exception_3,io_writeBackStage_inst_1_ex_exception_2,
    io_writeBackStage_inst_1_ex_exception_1,io_writeBackStage_inst_1_ex_exception_0}; // @[playground/src/defines/Util.scala 8:18]
  wire [15:0] _io_regfile_1_wen_T_9 = {io_writeBackStage_inst_1_ex_exception_15,1'h0,
    io_writeBackStage_inst_1_ex_exception_13,io_writeBackStage_inst_1_ex_exception_12,
    io_writeBackStage_inst_1_ex_exception_11,1'h0,io_writeBackStage_inst_1_ex_exception_9,
    io_writeBackStage_inst_1_ex_exception_8,io_regfile_1_wen_lo_2}; // @[playground/src/defines/Util.scala 8:18]
  wire [5:0] io_regfile_1_wen_lo_3 = {io_writeBackStage_inst_1_ex_interrupt_5,io_writeBackStage_inst_1_ex_interrupt_4,
    io_writeBackStage_inst_1_ex_interrupt_3,io_writeBackStage_inst_1_ex_interrupt_2,
    io_writeBackStage_inst_1_ex_interrupt_1,io_writeBackStage_inst_1_ex_interrupt_0}; // @[playground/src/defines/Util.scala 8:45]
  wire [11:0] _io_regfile_1_wen_T_11 = {io_writeBackStage_inst_1_ex_interrupt_11,
    io_writeBackStage_inst_1_ex_interrupt_10,io_writeBackStage_inst_1_ex_interrupt_9,
    io_writeBackStage_inst_1_ex_interrupt_8,io_writeBackStage_inst_1_ex_interrupt_7,
    io_writeBackStage_inst_1_ex_interrupt_6,io_regfile_1_wen_lo_3}; // @[playground/src/defines/Util.scala 8:45]
  wire  _io_regfile_1_wen_T_13 = |_io_regfile_1_wen_T_9 | |_io_regfile_1_wen_T_11; // @[playground/src/defines/Util.scala 8:29]
  wire  _io_regfile_1_wen_T_14 = ~_io_regfile_1_wen_T_13; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 29:7]
  wire [63:0] _GEN_1 = 3'h1 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_1 :
    io_writeBackStage_inst_0_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_2 = 3'h2 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_2 : _GEN_1; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_3 = 3'h3 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_3 : _GEN_2; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_4 = 3'h4 == io_writeBackStage_inst_0_info_fusel ? 64'h0 : _GEN_3; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_7 = 3'h1 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_1 :
    io_writeBackStage_inst_1_rd_info_wdata_0; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_8 = 3'h2 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_2 : _GEN_7; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_9 = 3'h3 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_3 : _GEN_8; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire [63:0] _GEN_10 = 3'h4 == io_writeBackStage_inst_1_info_fusel ? 64'h0 : _GEN_9; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  wire  _io_debug_wb_pc_T_2 = io_writeBackStage_inst_1_info_valid & io_ctrl_allow_to_go; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 54:48]
  wire  _io_debug_wb_pc_T_3 = ~(io_writeBackStage_inst_1_info_valid & io_ctrl_allow_to_go); // @[playground/src/pipeline/writeback/WriteBackUnit.scala 54:9]
  wire [63:0] _io_debug_wb_pc_T_4 = _io_debug_wb_pc_T_3 ? 64'h0 : io_writeBackStage_inst_1_pc; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 53:10]
  wire  _io_debug_wb_rf_wen_T_2 = io_writeBackStage_inst_0_info_valid & io_ctrl_allow_to_go; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 61:44]
  assign io_regfile_0_wen = _io_regfile_0_wen_T_1 & _io_regfile_0_wen_T_7; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 21:27]
  assign io_regfile_0_waddr = io_writeBackStage_inst_0_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 32:25]
  assign io_regfile_0_wdata = 3'h5 == io_writeBackStage_inst_0_info_fusel ? io_writeBackStage_inst_0_rd_info_wdata_5 :
    _GEN_4; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  assign io_regfile_1_wen = _io_regfile_1_wen_T_8 & _io_regfile_1_wen_T_14; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 28:50]
  assign io_regfile_1_waddr = io_writeBackStage_inst_1_info_reg_waddr; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 32:25]
  assign io_regfile_1_wdata = 3'h5 == io_writeBackStage_inst_1_info_fusel ? io_writeBackStage_inst_1_rd_info_wdata_5 :
    _GEN_10; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 33:{25,25}]
  assign io_debug_wb_pc = clock ? io_writeBackStage_inst_0_pc : _io_debug_wb_pc_T_4; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 50:26]
  assign io_debug_wb_rf_wen = clock ? _io_debug_wb_rf_wen_T_2 : _io_debug_wb_pc_T_2; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 59:30]
  assign io_debug_wb_rf_wnum = clock ? io_regfile_0_waddr : io_regfile_1_waddr; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 64:31]
  assign io_debug_wb_rf_wdata = clock ? io_regfile_0_wdata : io_regfile_1_wdata; // @[playground/src/pipeline/writeback/WriteBackUnit.scala 69:32]
endmodule
module Tlb(
  input         clock,
  input         reset,
  input         io_icache_en, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [63:0] io_icache_vaddr, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_icache_complete_single_request, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_icache_uncached, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_icache_hit, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [19:0] io_icache_ptag, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [31:0] io_icache_paddr, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_icache_page_fault, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_en, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [63:0] io_dcache_vaddr, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_complete_single_request, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_dcache_uncached, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_dcache_hit, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [19:0] io_dcache_ptag, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [31:0] io_dcache_paddr, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_dcache_page_fault, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [1:0]  io_dcache_access_type, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_vpn_ready, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output        io_dcache_ptw_vpn_valid, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [26:0] io_dcache_ptw_vpn_bits, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [1:0]  io_dcache_ptw_access_type, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_valid, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_page_fault, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [19:0] io_dcache_ptw_pte_bits_entry_ppn, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_d, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_g, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_u, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_x, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_w, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_r, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_dcache_ptw_pte_bits_entry_flag_v, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [17:0] io_dcache_ptw_pte_bits_rmask, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [63:0] io_dcache_csr_satp, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [63:0] io_dcache_csr_mstatus, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [1:0]  io_dcache_csr_imode, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  output [1:0]  io_dcache_csr_dmode, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [63:0] io_csr_satp, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [63:0] io_csr_mstatus, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [1:0]  io_csr_imode, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [1:0]  io_csr_dmode, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input         io_sfence_vma_valid, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [63:0] io_sfence_vma_src_info_src1_data, // @[playground/src/cache/mmu/Tlb.scala 51:14]
  input  [63:0] io_sfence_vma_src_info_src2_data // @[playground/src/cache/mmu/Tlb.scala 51:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] satp_asid = io_csr_satp[59:44]; // @[playground/src/cache/mmu/Tlb.scala 58:37]
  wire [3:0] satp_mode = io_csr_satp[63:60]; // @[playground/src/cache/mmu/Tlb.scala 58:37]
  wire  mstatus_sum = io_csr_mstatus[18]; // @[playground/src/cache/mmu/Tlb.scala 59:40]
  wire  mstatus_mxr = io_csr_mstatus[19]; // @[playground/src/cache/mmu/Tlb.scala 59:40]
  wire  _ivm_enabled_T = satp_mode == 4'h8; // @[playground/src/cache/mmu/Tlb.scala 72:32]
  wire  ivm_enabled = satp_mode == 4'h8 & io_csr_imode < 2'h3; // @[playground/src/cache/mmu/Tlb.scala 72:41]
  wire  dvm_enabled = _ivm_enabled_T & io_csr_dmode < 2'h3; // @[playground/src/cache/mmu/Tlb.scala 73:41]
  reg [26:0] itlb_vpn; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg [15:0] itlb_asid; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg  itlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg  itlb_flag_u; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg  itlb_flag_x; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg  itlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg [19:0] itlb_ppn; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg [17:0] itlb_rmask; // @[playground/src/cache/mmu/Tlb.scala 75:22]
  reg [26:0] dtlb_vpn; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg [15:0] dtlb_asid; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_d; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_u; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_x; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_w; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_r; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg  dtlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg [19:0] dtlb_ppn; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg [17:0] dtlb_rmask; // @[playground/src/cache/mmu/Tlb.scala 76:22]
  reg [26:0] tlbl2_0_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_0_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_0_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_0_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_1_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_1_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_1_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_1_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_1_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_2_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_2_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_2_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_2_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_2_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_3_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_3_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_3_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_3_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_3_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_4_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_4_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_4_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_4_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_4_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_5_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_5_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_5_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_5_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_5_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_6_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_6_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_6_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_6_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_6_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_7_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_7_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_7_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_7_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_7_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_8_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_8_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_8_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_8_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_8_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_9_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_9_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_9_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_9_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_9_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_10_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_10_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_10_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_10_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_10_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_11_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_11_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_11_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_11_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_11_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_12_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_12_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_12_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_12_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_12_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_13_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_13_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_13_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_13_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_13_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_14_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_14_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_14_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_14_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_14_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [26:0] tlbl2_15_vpn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [15:0] tlbl2_15_asid; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_d; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_g; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_u; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_x; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_w; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_r; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg  tlbl2_15_flag_v; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [19:0] tlbl2_15_ppn; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  reg [17:0] tlbl2_15_rmask; // @[playground/src/cache/mmu/Tlb.scala 77:22]
  wire [26:0] ivpn = io_icache_vaddr[38:12]; // @[playground/src/cache/mmu/Tlb.scala 79:29]
  wire [26:0] dvpn = io_dcache_vaddr[38:12]; // @[playground/src/cache/mmu/Tlb.scala 80:29]
  wire [26:0] itlbl1_hit_fullmask = {9'h1ff,itlb_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _itlbl1_hit_T = ivpn & itlbl1_hit_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _itlbl1_hit_T_1 = itlb_vpn & itlbl1_hit_fullmask; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _itlbl1_hit_T_2 = _itlbl1_hit_T == _itlbl1_hit_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _itlbl1_hit_T_4 = itlb_asid == satp_asid | itlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 84:30]
  wire  _itlbl1_hit_T_5 = _itlbl1_hit_T_2 & _itlbl1_hit_T_4; // @[playground/src/cache/mmu/Tlb.scala 83:54]
  wire  itlbl1_hit = _itlbl1_hit_T_5 & itlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 84:46]
  wire [26:0] dtlbl1_hit_fullmask = {9'h1ff,dtlb_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _dtlbl1_hit_T = dvpn & dtlbl1_hit_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _dtlbl1_hit_T_1 = dtlb_vpn & dtlbl1_hit_fullmask; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _dtlbl1_hit_T_2 = _dtlbl1_hit_T == _dtlbl1_hit_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dtlbl1_hit_T_4 = dtlb_asid == satp_asid | dtlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 87:30]
  wire  _dtlbl1_hit_T_5 = _dtlbl1_hit_T_2 & _dtlbl1_hit_T_4; // @[playground/src/cache/mmu/Tlb.scala 86:54]
  wire  dtlbl1_hit = _dtlbl1_hit_T_5 & dtlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 87:46]
  wire [26:0] il2_hit_vec_fullmask = {9'h1ff,tlbl2_0_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T = ivpn & il2_hit_vec_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_1 = tlbl2_0_vpn & il2_hit_vec_fullmask; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_2 = _il2_hit_vec_T == _il2_hit_vec_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_4 = tlbl2_0_asid == satp_asid | tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_5 = _il2_hit_vec_T_2 & _il2_hit_vec_T_4; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_0 = _il2_hit_vec_T_5 & tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_1 = {9'h1ff,tlbl2_1_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_7 = ivpn & il2_hit_vec_fullmask_1; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_8 = tlbl2_1_vpn & il2_hit_vec_fullmask_1; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_9 = _il2_hit_vec_T_7 == _il2_hit_vec_T_8; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_11 = tlbl2_1_asid == satp_asid | tlbl2_1_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_12 = _il2_hit_vec_T_9 & _il2_hit_vec_T_11; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_1 = _il2_hit_vec_T_12 & tlbl2_1_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_2 = {9'h1ff,tlbl2_2_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_14 = ivpn & il2_hit_vec_fullmask_2; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_15 = tlbl2_2_vpn & il2_hit_vec_fullmask_2; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_16 = _il2_hit_vec_T_14 == _il2_hit_vec_T_15; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_18 = tlbl2_2_asid == satp_asid | tlbl2_2_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_19 = _il2_hit_vec_T_16 & _il2_hit_vec_T_18; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_2 = _il2_hit_vec_T_19 & tlbl2_2_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_3 = {9'h1ff,tlbl2_3_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_21 = ivpn & il2_hit_vec_fullmask_3; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_22 = tlbl2_3_vpn & il2_hit_vec_fullmask_3; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_23 = _il2_hit_vec_T_21 == _il2_hit_vec_T_22; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_25 = tlbl2_3_asid == satp_asid | tlbl2_3_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_26 = _il2_hit_vec_T_23 & _il2_hit_vec_T_25; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_3 = _il2_hit_vec_T_26 & tlbl2_3_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_4 = {9'h1ff,tlbl2_4_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_28 = ivpn & il2_hit_vec_fullmask_4; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_29 = tlbl2_4_vpn & il2_hit_vec_fullmask_4; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_30 = _il2_hit_vec_T_28 == _il2_hit_vec_T_29; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_32 = tlbl2_4_asid == satp_asid | tlbl2_4_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_33 = _il2_hit_vec_T_30 & _il2_hit_vec_T_32; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_4 = _il2_hit_vec_T_33 & tlbl2_4_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_5 = {9'h1ff,tlbl2_5_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_35 = ivpn & il2_hit_vec_fullmask_5; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_36 = tlbl2_5_vpn & il2_hit_vec_fullmask_5; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_37 = _il2_hit_vec_T_35 == _il2_hit_vec_T_36; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_39 = tlbl2_5_asid == satp_asid | tlbl2_5_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_40 = _il2_hit_vec_T_37 & _il2_hit_vec_T_39; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_5 = _il2_hit_vec_T_40 & tlbl2_5_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_6 = {9'h1ff,tlbl2_6_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_42 = ivpn & il2_hit_vec_fullmask_6; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_43 = tlbl2_6_vpn & il2_hit_vec_fullmask_6; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_44 = _il2_hit_vec_T_42 == _il2_hit_vec_T_43; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_46 = tlbl2_6_asid == satp_asid | tlbl2_6_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_47 = _il2_hit_vec_T_44 & _il2_hit_vec_T_46; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_6 = _il2_hit_vec_T_47 & tlbl2_6_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_7 = {9'h1ff,tlbl2_7_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_49 = ivpn & il2_hit_vec_fullmask_7; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_50 = tlbl2_7_vpn & il2_hit_vec_fullmask_7; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_51 = _il2_hit_vec_T_49 == _il2_hit_vec_T_50; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_53 = tlbl2_7_asid == satp_asid | tlbl2_7_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_54 = _il2_hit_vec_T_51 & _il2_hit_vec_T_53; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_7 = _il2_hit_vec_T_54 & tlbl2_7_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_8 = {9'h1ff,tlbl2_8_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_56 = ivpn & il2_hit_vec_fullmask_8; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_57 = tlbl2_8_vpn & il2_hit_vec_fullmask_8; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_58 = _il2_hit_vec_T_56 == _il2_hit_vec_T_57; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_60 = tlbl2_8_asid == satp_asid | tlbl2_8_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_61 = _il2_hit_vec_T_58 & _il2_hit_vec_T_60; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_8 = _il2_hit_vec_T_61 & tlbl2_8_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_9 = {9'h1ff,tlbl2_9_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_63 = ivpn & il2_hit_vec_fullmask_9; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_64 = tlbl2_9_vpn & il2_hit_vec_fullmask_9; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_65 = _il2_hit_vec_T_63 == _il2_hit_vec_T_64; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_67 = tlbl2_9_asid == satp_asid | tlbl2_9_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_68 = _il2_hit_vec_T_65 & _il2_hit_vec_T_67; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_9 = _il2_hit_vec_T_68 & tlbl2_9_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_10 = {9'h1ff,tlbl2_10_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_70 = ivpn & il2_hit_vec_fullmask_10; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_71 = tlbl2_10_vpn & il2_hit_vec_fullmask_10; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_72 = _il2_hit_vec_T_70 == _il2_hit_vec_T_71; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_74 = tlbl2_10_asid == satp_asid | tlbl2_10_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_75 = _il2_hit_vec_T_72 & _il2_hit_vec_T_74; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_10 = _il2_hit_vec_T_75 & tlbl2_10_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_11 = {9'h1ff,tlbl2_11_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_77 = ivpn & il2_hit_vec_fullmask_11; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_78 = tlbl2_11_vpn & il2_hit_vec_fullmask_11; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_79 = _il2_hit_vec_T_77 == _il2_hit_vec_T_78; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_81 = tlbl2_11_asid == satp_asid | tlbl2_11_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_82 = _il2_hit_vec_T_79 & _il2_hit_vec_T_81; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_11 = _il2_hit_vec_T_82 & tlbl2_11_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_12 = {9'h1ff,tlbl2_12_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_84 = ivpn & il2_hit_vec_fullmask_12; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_85 = tlbl2_12_vpn & il2_hit_vec_fullmask_12; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_86 = _il2_hit_vec_T_84 == _il2_hit_vec_T_85; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_88 = tlbl2_12_asid == satp_asid | tlbl2_12_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_89 = _il2_hit_vec_T_86 & _il2_hit_vec_T_88; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_12 = _il2_hit_vec_T_89 & tlbl2_12_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_13 = {9'h1ff,tlbl2_13_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_91 = ivpn & il2_hit_vec_fullmask_13; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_92 = tlbl2_13_vpn & il2_hit_vec_fullmask_13; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_93 = _il2_hit_vec_T_91 == _il2_hit_vec_T_92; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_95 = tlbl2_13_asid == satp_asid | tlbl2_13_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_96 = _il2_hit_vec_T_93 & _il2_hit_vec_T_95; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_13 = _il2_hit_vec_T_96 & tlbl2_13_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_14 = {9'h1ff,tlbl2_14_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_98 = ivpn & il2_hit_vec_fullmask_14; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_99 = tlbl2_14_vpn & il2_hit_vec_fullmask_14; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_100 = _il2_hit_vec_T_98 == _il2_hit_vec_T_99; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_102 = tlbl2_14_asid == satp_asid | tlbl2_14_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_103 = _il2_hit_vec_T_100 & _il2_hit_vec_T_102; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_14 = _il2_hit_vec_T_103 & tlbl2_14_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] il2_hit_vec_fullmask_15 = {9'h1ff,tlbl2_15_rmask}; // @[playground/src/defines/TlbBundles.scala 36:23]
  wire [26:0] _il2_hit_vec_T_105 = ivpn & il2_hit_vec_fullmask_15; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _il2_hit_vec_T_106 = tlbl2_15_vpn & il2_hit_vec_fullmask_15; // @[playground/src/defines/TlbBundles.scala 37:34]
  wire  _il2_hit_vec_T_107 = _il2_hit_vec_T_105 == _il2_hit_vec_T_106; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _il2_hit_vec_T_109 = tlbl2_15_asid == satp_asid | tlbl2_15_flag_g; // @[playground/src/cache/mmu/Tlb.scala 93:33]
  wire  _il2_hit_vec_T_110 = _il2_hit_vec_T_107 & _il2_hit_vec_T_109; // @[playground/src/cache/mmu/Tlb.scala 92:39]
  wire  il2_hit_vec_15 = _il2_hit_vec_T_110 & tlbl2_15_flag_v; // @[playground/src/cache/mmu/Tlb.scala 93:48]
  wire [26:0] _dl2_hit_vec_T = dvpn & il2_hit_vec_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_2 = _dl2_hit_vec_T == _il2_hit_vec_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_5 = _dl2_hit_vec_T_2 & _il2_hit_vec_T_4; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_0 = _dl2_hit_vec_T_5 & tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_7 = dvpn & il2_hit_vec_fullmask_1; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_9 = _dl2_hit_vec_T_7 == _il2_hit_vec_T_8; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_12 = _dl2_hit_vec_T_9 & _il2_hit_vec_T_11; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_1 = _dl2_hit_vec_T_12 & tlbl2_1_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_14 = dvpn & il2_hit_vec_fullmask_2; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_16 = _dl2_hit_vec_T_14 == _il2_hit_vec_T_15; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_19 = _dl2_hit_vec_T_16 & _il2_hit_vec_T_18; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_2 = _dl2_hit_vec_T_19 & tlbl2_2_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_21 = dvpn & il2_hit_vec_fullmask_3; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_23 = _dl2_hit_vec_T_21 == _il2_hit_vec_T_22; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_26 = _dl2_hit_vec_T_23 & _il2_hit_vec_T_25; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_3 = _dl2_hit_vec_T_26 & tlbl2_3_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_28 = dvpn & il2_hit_vec_fullmask_4; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_30 = _dl2_hit_vec_T_28 == _il2_hit_vec_T_29; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_33 = _dl2_hit_vec_T_30 & _il2_hit_vec_T_32; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_4 = _dl2_hit_vec_T_33 & tlbl2_4_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_35 = dvpn & il2_hit_vec_fullmask_5; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_37 = _dl2_hit_vec_T_35 == _il2_hit_vec_T_36; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_40 = _dl2_hit_vec_T_37 & _il2_hit_vec_T_39; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_5 = _dl2_hit_vec_T_40 & tlbl2_5_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_42 = dvpn & il2_hit_vec_fullmask_6; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_44 = _dl2_hit_vec_T_42 == _il2_hit_vec_T_43; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_47 = _dl2_hit_vec_T_44 & _il2_hit_vec_T_46; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_6 = _dl2_hit_vec_T_47 & tlbl2_6_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_49 = dvpn & il2_hit_vec_fullmask_7; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_51 = _dl2_hit_vec_T_49 == _il2_hit_vec_T_50; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_54 = _dl2_hit_vec_T_51 & _il2_hit_vec_T_53; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_7 = _dl2_hit_vec_T_54 & tlbl2_7_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_56 = dvpn & il2_hit_vec_fullmask_8; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_58 = _dl2_hit_vec_T_56 == _il2_hit_vec_T_57; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_61 = _dl2_hit_vec_T_58 & _il2_hit_vec_T_60; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_8 = _dl2_hit_vec_T_61 & tlbl2_8_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_63 = dvpn & il2_hit_vec_fullmask_9; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_65 = _dl2_hit_vec_T_63 == _il2_hit_vec_T_64; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_68 = _dl2_hit_vec_T_65 & _il2_hit_vec_T_67; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_9 = _dl2_hit_vec_T_68 & tlbl2_9_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_70 = dvpn & il2_hit_vec_fullmask_10; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_72 = _dl2_hit_vec_T_70 == _il2_hit_vec_T_71; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_75 = _dl2_hit_vec_T_72 & _il2_hit_vec_T_74; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_10 = _dl2_hit_vec_T_75 & tlbl2_10_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_77 = dvpn & il2_hit_vec_fullmask_11; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_79 = _dl2_hit_vec_T_77 == _il2_hit_vec_T_78; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_82 = _dl2_hit_vec_T_79 & _il2_hit_vec_T_81; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_11 = _dl2_hit_vec_T_82 & tlbl2_11_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_84 = dvpn & il2_hit_vec_fullmask_12; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_86 = _dl2_hit_vec_T_84 == _il2_hit_vec_T_85; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_89 = _dl2_hit_vec_T_86 & _il2_hit_vec_T_88; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_12 = _dl2_hit_vec_T_89 & tlbl2_12_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_91 = dvpn & il2_hit_vec_fullmask_13; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_93 = _dl2_hit_vec_T_91 == _il2_hit_vec_T_92; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_96 = _dl2_hit_vec_T_93 & _il2_hit_vec_T_95; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_13 = _dl2_hit_vec_T_96 & tlbl2_13_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_98 = dvpn & il2_hit_vec_fullmask_14; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_100 = _dl2_hit_vec_T_98 == _il2_hit_vec_T_99; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_103 = _dl2_hit_vec_T_100 & _il2_hit_vec_T_102; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_14 = _dl2_hit_vec_T_103 & tlbl2_14_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  wire [26:0] _dl2_hit_vec_T_105 = dvpn & il2_hit_vec_fullmask_15; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _dl2_hit_vec_T_107 = _dl2_hit_vec_T_105 == _il2_hit_vec_T_106; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _dl2_hit_vec_T_110 = _dl2_hit_vec_T_107 & _il2_hit_vec_T_109; // @[playground/src/cache/mmu/Tlb.scala 99:39]
  wire  dl2_hit_vec_15 = _dl2_hit_vec_T_110 & tlbl2_15_flag_v; // @[playground/src/cache/mmu/Tlb.scala 100:48]
  reg [1:0] immu_state; // @[playground/src/cache/mmu/Tlb.scala 106:76]
  reg [1:0] dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 107:76]
  reg [3:0] replace_index_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  ipage_fault; // @[playground/src/cache/mmu/Tlb.scala 112:30]
  reg  dpage_fault; // @[playground/src/cache/mmu/Tlb.scala 113:30]
  reg  ar_sel_lock; // @[playground/src/cache/mmu/Tlb.scala 120:28]
  reg  ar_sel_val; // @[playground/src/cache/mmu/Tlb.scala 121:28]
  wire [7:0] lo_1 = {dl2_hit_vec_7,dl2_hit_vec_6,dl2_hit_vec_5,dl2_hit_vec_4,dl2_hit_vec_3,dl2_hit_vec_2,dl2_hit_vec_1,
    dl2_hit_vec_0}; // @[playground/src/cache/mmu/Tlb.scala 320:24]
  wire [15:0] _T_40 = {dl2_hit_vec_15,dl2_hit_vec_14,dl2_hit_vec_13,dl2_hit_vec_12,dl2_hit_vec_11,dl2_hit_vec_10,
    dl2_hit_vec_9,dl2_hit_vec_8,lo_1}; // @[playground/src/cache/mmu/Tlb.scala 320:24]
  wire  _GEN_1958 = |_T_40 ? 1'h0 : 1'h1; // @[playground/src/cache/mmu/Tlb.scala 118:25 320:36 324:20]
  wire  _GEN_3000 = 2'h1 == dmmu_state ? _GEN_1958 : 2'h2 == dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  req_ptw_1 = 2'h0 == dmmu_state ? 1'h0 : _GEN_3000; // @[playground/src/cache/mmu/Tlb.scala 266:22 118:25]
  wire [7:0] lo = {il2_hit_vec_7,il2_hit_vec_6,il2_hit_vec_5,il2_hit_vec_4,il2_hit_vec_3,il2_hit_vec_2,il2_hit_vec_1,
    il2_hit_vec_0}; // @[playground/src/cache/mmu/Tlb.scala 220:24]
  wire [15:0] _T_9 = {il2_hit_vec_15,il2_hit_vec_14,il2_hit_vec_13,il2_hit_vec_12,il2_hit_vec_11,il2_hit_vec_10,
    il2_hit_vec_9,il2_hit_vec_8,lo}; // @[playground/src/cache/mmu/Tlb.scala 220:24]
  wire  _GEN_235 = |_T_9 ? 1'h0 : 1'h1; // @[playground/src/cache/mmu/Tlb.scala 118:25 220:36 224:20]
  wire  _GEN_1279 = 2'h1 == immu_state ? _GEN_235 : 2'h2 == immu_state; // @[playground/src/cache/mmu/Tlb.scala 193:22]
  wire  req_ptw_0 = 2'h0 == immu_state ? 1'h0 : _GEN_1279; // @[playground/src/cache/mmu/Tlb.scala 193:22 118:25]
  wire  choose_icache = ar_sel_lock ? ar_sel_val : req_ptw_0 & ~req_ptw_1; // @[playground/src/cache/mmu/Tlb.scala 123:26]
  wire  _T_4 = ~mstatus_sum; // @[playground/src/cache/mmu/Tlb.scala 151:33]
  wire  _T_5 = itlb_flag_u & ~mstatus_sum; // @[playground/src/cache/mmu/Tlb.scala 151:26]
  wire [1:0] _GEN_5 = itlb_flag_u & ~mstatus_sum ? 2'h3 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 151:42 153:23 106:76]
  wire  _GEN_6 = itlb_flag_u & ~mstatus_sum ? 1'h0 : 1'h1; // @[playground/src/cache/mmu/Tlb.scala 151:42 155:25 207:25]
  wire  _T_7 = ~itlb_flag_u; // @[playground/src/cache/mmu/Tlb.scala 159:14]
  wire [1:0] _GEN_8 = ~itlb_flag_u ? 2'h3 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 159:28 161:23 106:76]
  wire  _GEN_9 = ~itlb_flag_u ? 1'h0 : 1'h1; // @[playground/src/cache/mmu/Tlb.scala 159:28 163:25 207:25]
  wire  _GEN_10 = 2'h0 == io_csr_imode & _T_7; // @[playground/src/cache/mmu/Tlb.scala 149:19 197:23]
  wire [1:0] _GEN_11 = 2'h0 == io_csr_imode ? _GEN_8 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 149:19 106:76]
  wire  _GEN_12 = 2'h0 == io_csr_imode & _GEN_9; // @[playground/src/cache/mmu/Tlb.scala 149:19 207:25]
  wire  _GEN_13 = 2'h1 == io_csr_imode ? _T_5 : _GEN_10; // @[playground/src/cache/mmu/Tlb.scala 149:19]
  wire [1:0] _GEN_14 = 2'h1 == io_csr_imode ? _GEN_5 : _GEN_11; // @[playground/src/cache/mmu/Tlb.scala 149:19]
  wire  _GEN_15 = 2'h1 == io_csr_imode ? _GEN_6 : _GEN_12; // @[playground/src/cache/mmu/Tlb.scala 149:19]
  wire  _GEN_16 = ~itlb_flag_x | _GEN_13; // @[playground/src/cache/mmu/Tlb.scala 208:30 209:25]
  wire [1:0] _GEN_17 = ~itlb_flag_x ? 2'h3 : _GEN_14; // @[playground/src/cache/mmu/Tlb.scala 208:30 210:25]
  wire  _GEN_18 = ~itlb_flag_x ? 1'h0 : _GEN_15; // @[playground/src/cache/mmu/Tlb.scala 207:25 208:30]
  wire  _GEN_19 = itlbl1_hit & _GEN_18; // @[playground/src/cache/mmu/Tlb.scala 134:26 201:32]
  wire  _GEN_20 = itlbl1_hit & _GEN_16; // @[playground/src/cache/mmu/Tlb.scala 197:23 201:32]
  wire [1:0] _GEN_21 = itlbl1_hit ? _GEN_17 : 2'h1; // @[playground/src/cache/mmu/Tlb.scala 201:32 215:22]
  wire  _GEN_22 = ~ivm_enabled | _GEN_19; // @[playground/src/cache/mmu/Tlb.scala 199:28 200:25]
  wire  _GEN_27 = io_icache_en & _GEN_22; // @[playground/src/cache/mmu/Tlb.scala 134:26 195:26]
  wire [3:0] _itlb_T = il2_hit_vec_14 ? 4'he : 4'hf; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_1 = il2_hit_vec_13 ? 4'hd : _itlb_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_2 = il2_hit_vec_12 ? 4'hc : _itlb_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_3 = il2_hit_vec_11 ? 4'hb : _itlb_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_4 = il2_hit_vec_10 ? 4'ha : _itlb_T_3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_5 = il2_hit_vec_9 ? 4'h9 : _itlb_T_4; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_6 = il2_hit_vec_8 ? 4'h8 : _itlb_T_5; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_7 = il2_hit_vec_7 ? 4'h7 : _itlb_T_6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_8 = il2_hit_vec_6 ? 4'h6 : _itlb_T_7; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_9 = il2_hit_vec_5 ? 4'h5 : _itlb_T_8; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_10 = il2_hit_vec_4 ? 4'h4 : _itlb_T_9; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_11 = il2_hit_vec_3 ? 4'h3 : _itlb_T_10; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_12 = il2_hit_vec_2 ? 4'h2 : _itlb_T_11; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_13 = il2_hit_vec_1 ? 4'h1 : _itlb_T_12; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _itlb_T_14 = il2_hit_vec_0 ? 4'h0 : _itlb_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [26:0] _GEN_30 = 4'h1 == _itlb_T_14 ? tlbl2_1_vpn : tlbl2_0_vpn; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_31 = 4'h2 == _itlb_T_14 ? tlbl2_2_vpn : _GEN_30; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_32 = 4'h3 == _itlb_T_14 ? tlbl2_3_vpn : _GEN_31; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_33 = 4'h4 == _itlb_T_14 ? tlbl2_4_vpn : _GEN_32; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_34 = 4'h5 == _itlb_T_14 ? tlbl2_5_vpn : _GEN_33; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_35 = 4'h6 == _itlb_T_14 ? tlbl2_6_vpn : _GEN_34; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_36 = 4'h7 == _itlb_T_14 ? tlbl2_7_vpn : _GEN_35; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_37 = 4'h8 == _itlb_T_14 ? tlbl2_8_vpn : _GEN_36; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_38 = 4'h9 == _itlb_T_14 ? tlbl2_9_vpn : _GEN_37; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_39 = 4'ha == _itlb_T_14 ? tlbl2_10_vpn : _GEN_38; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_40 = 4'hb == _itlb_T_14 ? tlbl2_11_vpn : _GEN_39; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_41 = 4'hc == _itlb_T_14 ? tlbl2_12_vpn : _GEN_40; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_42 = 4'hd == _itlb_T_14 ? tlbl2_13_vpn : _GEN_41; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_43 = 4'he == _itlb_T_14 ? tlbl2_14_vpn : _GEN_42; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [26:0] _GEN_44 = 4'hf == _itlb_T_14 ? tlbl2_15_vpn : _GEN_43; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_46 = 4'h1 == _itlb_T_14 ? tlbl2_1_asid : tlbl2_0_asid; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_47 = 4'h2 == _itlb_T_14 ? tlbl2_2_asid : _GEN_46; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_48 = 4'h3 == _itlb_T_14 ? tlbl2_3_asid : _GEN_47; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_49 = 4'h4 == _itlb_T_14 ? tlbl2_4_asid : _GEN_48; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_50 = 4'h5 == _itlb_T_14 ? tlbl2_5_asid : _GEN_49; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_51 = 4'h6 == _itlb_T_14 ? tlbl2_6_asid : _GEN_50; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_52 = 4'h7 == _itlb_T_14 ? tlbl2_7_asid : _GEN_51; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_53 = 4'h8 == _itlb_T_14 ? tlbl2_8_asid : _GEN_52; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_54 = 4'h9 == _itlb_T_14 ? tlbl2_9_asid : _GEN_53; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_55 = 4'ha == _itlb_T_14 ? tlbl2_10_asid : _GEN_54; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_56 = 4'hb == _itlb_T_14 ? tlbl2_11_asid : _GEN_55; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_57 = 4'hc == _itlb_T_14 ? tlbl2_12_asid : _GEN_56; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_58 = 4'hd == _itlb_T_14 ? tlbl2_13_asid : _GEN_57; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_59 = 4'he == _itlb_T_14 ? tlbl2_14_asid : _GEN_58; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [15:0] _GEN_60 = 4'hf == _itlb_T_14 ? tlbl2_15_asid : _GEN_59; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_94 = 4'h1 == _itlb_T_14 ? tlbl2_1_flag_g : tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_95 = 4'h2 == _itlb_T_14 ? tlbl2_2_flag_g : _GEN_94; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_96 = 4'h3 == _itlb_T_14 ? tlbl2_3_flag_g : _GEN_95; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_97 = 4'h4 == _itlb_T_14 ? tlbl2_4_flag_g : _GEN_96; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_98 = 4'h5 == _itlb_T_14 ? tlbl2_5_flag_g : _GEN_97; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_99 = 4'h6 == _itlb_T_14 ? tlbl2_6_flag_g : _GEN_98; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_100 = 4'h7 == _itlb_T_14 ? tlbl2_7_flag_g : _GEN_99; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_101 = 4'h8 == _itlb_T_14 ? tlbl2_8_flag_g : _GEN_100; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_102 = 4'h9 == _itlb_T_14 ? tlbl2_9_flag_g : _GEN_101; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_103 = 4'ha == _itlb_T_14 ? tlbl2_10_flag_g : _GEN_102; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_104 = 4'hb == _itlb_T_14 ? tlbl2_11_flag_g : _GEN_103; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_105 = 4'hc == _itlb_T_14 ? tlbl2_12_flag_g : _GEN_104; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_106 = 4'hd == _itlb_T_14 ? tlbl2_13_flag_g : _GEN_105; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_107 = 4'he == _itlb_T_14 ? tlbl2_14_flag_g : _GEN_106; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_108 = 4'hf == _itlb_T_14 ? tlbl2_15_flag_g : _GEN_107; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_110 = 4'h1 == _itlb_T_14 ? tlbl2_1_flag_u : tlbl2_0_flag_u; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_111 = 4'h2 == _itlb_T_14 ? tlbl2_2_flag_u : _GEN_110; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_112 = 4'h3 == _itlb_T_14 ? tlbl2_3_flag_u : _GEN_111; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_113 = 4'h4 == _itlb_T_14 ? tlbl2_4_flag_u : _GEN_112; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_114 = 4'h5 == _itlb_T_14 ? tlbl2_5_flag_u : _GEN_113; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_115 = 4'h6 == _itlb_T_14 ? tlbl2_6_flag_u : _GEN_114; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_116 = 4'h7 == _itlb_T_14 ? tlbl2_7_flag_u : _GEN_115; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_117 = 4'h8 == _itlb_T_14 ? tlbl2_8_flag_u : _GEN_116; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_118 = 4'h9 == _itlb_T_14 ? tlbl2_9_flag_u : _GEN_117; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_119 = 4'ha == _itlb_T_14 ? tlbl2_10_flag_u : _GEN_118; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_120 = 4'hb == _itlb_T_14 ? tlbl2_11_flag_u : _GEN_119; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_121 = 4'hc == _itlb_T_14 ? tlbl2_12_flag_u : _GEN_120; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_122 = 4'hd == _itlb_T_14 ? tlbl2_13_flag_u : _GEN_121; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_123 = 4'he == _itlb_T_14 ? tlbl2_14_flag_u : _GEN_122; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_124 = 4'hf == _itlb_T_14 ? tlbl2_15_flag_u : _GEN_123; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_126 = 4'h1 == _itlb_T_14 ? tlbl2_1_flag_x : tlbl2_0_flag_x; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_127 = 4'h2 == _itlb_T_14 ? tlbl2_2_flag_x : _GEN_126; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_128 = 4'h3 == _itlb_T_14 ? tlbl2_3_flag_x : _GEN_127; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_129 = 4'h4 == _itlb_T_14 ? tlbl2_4_flag_x : _GEN_128; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_130 = 4'h5 == _itlb_T_14 ? tlbl2_5_flag_x : _GEN_129; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_131 = 4'h6 == _itlb_T_14 ? tlbl2_6_flag_x : _GEN_130; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_132 = 4'h7 == _itlb_T_14 ? tlbl2_7_flag_x : _GEN_131; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_133 = 4'h8 == _itlb_T_14 ? tlbl2_8_flag_x : _GEN_132; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_134 = 4'h9 == _itlb_T_14 ? tlbl2_9_flag_x : _GEN_133; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_135 = 4'ha == _itlb_T_14 ? tlbl2_10_flag_x : _GEN_134; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_136 = 4'hb == _itlb_T_14 ? tlbl2_11_flag_x : _GEN_135; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_137 = 4'hc == _itlb_T_14 ? tlbl2_12_flag_x : _GEN_136; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_138 = 4'hd == _itlb_T_14 ? tlbl2_13_flag_x : _GEN_137; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_139 = 4'he == _itlb_T_14 ? tlbl2_14_flag_x : _GEN_138; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_140 = 4'hf == _itlb_T_14 ? tlbl2_15_flag_x : _GEN_139; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_174 = 4'h1 == _itlb_T_14 ? tlbl2_1_flag_v : tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_175 = 4'h2 == _itlb_T_14 ? tlbl2_2_flag_v : _GEN_174; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_176 = 4'h3 == _itlb_T_14 ? tlbl2_3_flag_v : _GEN_175; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_177 = 4'h4 == _itlb_T_14 ? tlbl2_4_flag_v : _GEN_176; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_178 = 4'h5 == _itlb_T_14 ? tlbl2_5_flag_v : _GEN_177; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_179 = 4'h6 == _itlb_T_14 ? tlbl2_6_flag_v : _GEN_178; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_180 = 4'h7 == _itlb_T_14 ? tlbl2_7_flag_v : _GEN_179; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_181 = 4'h8 == _itlb_T_14 ? tlbl2_8_flag_v : _GEN_180; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_182 = 4'h9 == _itlb_T_14 ? tlbl2_9_flag_v : _GEN_181; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_183 = 4'ha == _itlb_T_14 ? tlbl2_10_flag_v : _GEN_182; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_184 = 4'hb == _itlb_T_14 ? tlbl2_11_flag_v : _GEN_183; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_185 = 4'hc == _itlb_T_14 ? tlbl2_12_flag_v : _GEN_184; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_186 = 4'hd == _itlb_T_14 ? tlbl2_13_flag_v : _GEN_185; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_187 = 4'he == _itlb_T_14 ? tlbl2_14_flag_v : _GEN_186; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire  _GEN_188 = 4'hf == _itlb_T_14 ? tlbl2_15_flag_v : _GEN_187; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_190 = 4'h1 == _itlb_T_14 ? tlbl2_1_ppn : tlbl2_0_ppn; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_191 = 4'h2 == _itlb_T_14 ? tlbl2_2_ppn : _GEN_190; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_192 = 4'h3 == _itlb_T_14 ? tlbl2_3_ppn : _GEN_191; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_193 = 4'h4 == _itlb_T_14 ? tlbl2_4_ppn : _GEN_192; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_194 = 4'h5 == _itlb_T_14 ? tlbl2_5_ppn : _GEN_193; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_195 = 4'h6 == _itlb_T_14 ? tlbl2_6_ppn : _GEN_194; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_196 = 4'h7 == _itlb_T_14 ? tlbl2_7_ppn : _GEN_195; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_197 = 4'h8 == _itlb_T_14 ? tlbl2_8_ppn : _GEN_196; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_198 = 4'h9 == _itlb_T_14 ? tlbl2_9_ppn : _GEN_197; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_199 = 4'ha == _itlb_T_14 ? tlbl2_10_ppn : _GEN_198; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_200 = 4'hb == _itlb_T_14 ? tlbl2_11_ppn : _GEN_199; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_201 = 4'hc == _itlb_T_14 ? tlbl2_12_ppn : _GEN_200; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_202 = 4'hd == _itlb_T_14 ? tlbl2_13_ppn : _GEN_201; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_203 = 4'he == _itlb_T_14 ? tlbl2_14_ppn : _GEN_202; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [19:0] _GEN_204 = 4'hf == _itlb_T_14 ? tlbl2_15_ppn : _GEN_203; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_206 = 4'h1 == _itlb_T_14 ? tlbl2_1_rmask : tlbl2_0_rmask; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_207 = 4'h2 == _itlb_T_14 ? tlbl2_2_rmask : _GEN_206; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_208 = 4'h3 == _itlb_T_14 ? tlbl2_3_rmask : _GEN_207; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_209 = 4'h4 == _itlb_T_14 ? tlbl2_4_rmask : _GEN_208; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_210 = 4'h5 == _itlb_T_14 ? tlbl2_5_rmask : _GEN_209; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_211 = 4'h6 == _itlb_T_14 ? tlbl2_6_rmask : _GEN_210; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_212 = 4'h7 == _itlb_T_14 ? tlbl2_7_rmask : _GEN_211; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_213 = 4'h8 == _itlb_T_14 ? tlbl2_8_rmask : _GEN_212; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_214 = 4'h9 == _itlb_T_14 ? tlbl2_9_rmask : _GEN_213; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_215 = 4'ha == _itlb_T_14 ? tlbl2_10_rmask : _GEN_214; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_216 = 4'hb == _itlb_T_14 ? tlbl2_11_rmask : _GEN_215; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_217 = 4'hc == _itlb_T_14 ? tlbl2_12_rmask : _GEN_216; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_218 = 4'hd == _itlb_T_14 ? tlbl2_13_rmask : _GEN_217; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_219 = 4'he == _itlb_T_14 ? tlbl2_14_rmask : _GEN_218; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [17:0] _GEN_220 = 4'hf == _itlb_T_14 ? tlbl2_15_rmask : _GEN_219; // @[playground/src/cache/mmu/Tlb.scala 222:{20,20}]
  wire [1:0] _GEN_221 = choose_icache & io_dcache_ptw_vpn_ready ? 2'h2 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 225:56 226:22 106:76]
  wire  _GEN_232 = |_T_9 ? _GEN_188 : itlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 220:36 222:20 75:22]
  wire [26:0] _GEN_236 = 4'h0 == replace_index_value ? ivpn : tlbl2_0_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_237 = 4'h1 == replace_index_value ? ivpn : tlbl2_1_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_238 = 4'h2 == replace_index_value ? ivpn : tlbl2_2_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_239 = 4'h3 == replace_index_value ? ivpn : tlbl2_3_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_240 = 4'h4 == replace_index_value ? ivpn : tlbl2_4_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_241 = 4'h5 == replace_index_value ? ivpn : tlbl2_5_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_242 = 4'h6 == replace_index_value ? ivpn : tlbl2_6_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_243 = 4'h7 == replace_index_value ? ivpn : tlbl2_7_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_244 = 4'h8 == replace_index_value ? ivpn : tlbl2_8_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_245 = 4'h9 == replace_index_value ? ivpn : tlbl2_9_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_246 = 4'ha == replace_index_value ? ivpn : tlbl2_10_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_247 = 4'hb == replace_index_value ? ivpn : tlbl2_11_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_248 = 4'hc == replace_index_value ? ivpn : tlbl2_12_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_249 = 4'hd == replace_index_value ? ivpn : tlbl2_13_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_250 = 4'he == replace_index_value ? ivpn : tlbl2_14_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [26:0] _GEN_251 = 4'hf == replace_index_value ? ivpn : tlbl2_15_vpn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_252 = 4'h0 == replace_index_value ? satp_asid : tlbl2_0_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_253 = 4'h1 == replace_index_value ? satp_asid : tlbl2_1_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_254 = 4'h2 == replace_index_value ? satp_asid : tlbl2_2_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_255 = 4'h3 == replace_index_value ? satp_asid : tlbl2_3_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_256 = 4'h4 == replace_index_value ? satp_asid : tlbl2_4_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_257 = 4'h5 == replace_index_value ? satp_asid : tlbl2_5_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_258 = 4'h6 == replace_index_value ? satp_asid : tlbl2_6_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_259 = 4'h7 == replace_index_value ? satp_asid : tlbl2_7_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_260 = 4'h8 == replace_index_value ? satp_asid : tlbl2_8_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_261 = 4'h9 == replace_index_value ? satp_asid : tlbl2_9_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_262 = 4'ha == replace_index_value ? satp_asid : tlbl2_10_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_263 = 4'hb == replace_index_value ? satp_asid : tlbl2_11_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_264 = 4'hc == replace_index_value ? satp_asid : tlbl2_12_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_265 = 4'hd == replace_index_value ? satp_asid : tlbl2_13_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_266 = 4'he == replace_index_value ? satp_asid : tlbl2_14_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [15:0] _GEN_267 = 4'hf == replace_index_value ? satp_asid : tlbl2_15_asid; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_268 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_0_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_269 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_1_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_270 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_2_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_271 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_3_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_272 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_4_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_273 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_5_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_274 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_6_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_275 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_7_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_276 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_8_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_277 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_9_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_278 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_10_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_279 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_11_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_280 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_12_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_281 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_13_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_282 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_14_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_283 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : tlbl2_15_flag_d; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_300 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_301 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_1_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_302 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_2_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_303 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_3_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_304 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_4_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_305 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_5_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_306 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_6_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_307 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_7_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_308 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_8_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_309 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_9_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_310 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_10_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_311 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_11_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_312 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_12_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_313 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_13_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_314 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_14_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_315 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : tlbl2_15_flag_g; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_316 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_0_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_317 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_1_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_318 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_2_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_319 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_3_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_320 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_4_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_321 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_5_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_322 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_6_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_323 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_7_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_324 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_8_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_325 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_9_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_326 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_10_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_327 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_11_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_328 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_12_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_329 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_13_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_330 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_14_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_331 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : tlbl2_15_flag_u; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_332 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_0_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_333 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_1_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_334 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_2_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_335 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_3_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_336 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_4_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_337 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_5_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_338 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_6_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_339 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_7_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_340 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_8_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_341 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_9_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_342 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_10_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_343 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_11_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_344 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_12_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_345 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_13_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_346 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_14_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_347 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : tlbl2_15_flag_x; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_348 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_0_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_349 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_1_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_350 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_2_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_351 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_3_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_352 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_4_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_353 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_5_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_354 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_6_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_355 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_7_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_356 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_8_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_357 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_9_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_358 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_10_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_359 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_11_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_360 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_12_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_361 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_13_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_362 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_14_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_363 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : tlbl2_15_flag_w; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_364 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_0_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_365 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_1_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_366 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_2_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_367 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_3_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_368 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_4_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_369 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_5_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_370 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_6_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_371 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_7_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_372 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_8_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_373 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_9_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_374 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_10_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_375 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_11_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_376 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_12_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_377 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_13_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_378 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_14_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_379 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : tlbl2_15_flag_r; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_380 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_381 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_1_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_382 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_2_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_383 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_3_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_384 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_4_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_385 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_5_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_386 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_6_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_387 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_7_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_388 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_8_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_389 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_9_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_390 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_10_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_391 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_11_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_392 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_12_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_393 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_13_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_394 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_14_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire  _GEN_395 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : tlbl2_15_flag_v; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_396 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_0_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_397 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_1_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_398 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_2_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_399 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_3_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_400 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_4_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_401 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_5_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_402 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_6_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_403 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_7_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_404 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_8_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_405 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_9_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_406 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_10_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_407 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_11_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_408 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_12_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_409 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_13_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_410 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_14_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [19:0] _GEN_411 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : tlbl2_15_ppn; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_412 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_0_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_413 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_1_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_414 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_2_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_415 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_3_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_416 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_4_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_417 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_5_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_418 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_6_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_419 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_7_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_420 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_8_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_421 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_9_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_422 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_10_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_423 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_11_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_424 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_12_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_425 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_13_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_426 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_14_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [17:0] _GEN_427 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_rmask : tlbl2_15_rmask; // @[playground/src/cache/mmu/Tlb.scala 247:{38,38} 77:22]
  wire [3:0] _value_T_1 = replace_index_value + 4'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _GEN_428 = io_dcache_ptw_pte_bits_page_fault | ipage_fault; // @[playground/src/cache/mmu/Tlb.scala 236:55 237:23 112:30]
  wire [1:0] _GEN_429 = io_dcache_ptw_pte_bits_page_fault ? 2'h3 : 2'h0; // @[playground/src/cache/mmu/Tlb.scala 236:55 238:23 250:22]
  wire [26:0] _GEN_430 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_vpn : _GEN_236; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_431 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_vpn : _GEN_237; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_432 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_vpn : _GEN_238; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_433 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_vpn : _GEN_239; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_434 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_vpn : _GEN_240; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_435 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_vpn : _GEN_241; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_436 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_vpn : _GEN_242; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_437 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_vpn : _GEN_243; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_438 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_vpn : _GEN_244; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_439 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_vpn : _GEN_245; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_440 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_vpn : _GEN_246; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_441 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_vpn : _GEN_247; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_442 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_vpn : _GEN_248; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_443 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_vpn : _GEN_249; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_444 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_vpn : _GEN_250; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_445 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_vpn : _GEN_251; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_446 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_asid : _GEN_252; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_447 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_asid : _GEN_253; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_448 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_asid : _GEN_254; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_449 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_asid : _GEN_255; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_450 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_asid : _GEN_256; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_451 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_asid : _GEN_257; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_452 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_asid : _GEN_258; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_453 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_asid : _GEN_259; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_454 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_asid : _GEN_260; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_455 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_asid : _GEN_261; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_456 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_asid : _GEN_262; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_457 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_asid : _GEN_263; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_458 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_asid : _GEN_264; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_459 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_asid : _GEN_265; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_460 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_asid : _GEN_266; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [15:0] _GEN_461 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_asid : _GEN_267; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_462 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_d : _GEN_268; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_463 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_d : _GEN_269; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_464 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_d : _GEN_270; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_465 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_d : _GEN_271; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_466 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_d : _GEN_272; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_467 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_d : _GEN_273; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_468 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_d : _GEN_274; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_469 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_d : _GEN_275; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_470 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_d : _GEN_276; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_471 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_d : _GEN_277; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_472 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_d : _GEN_278; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_473 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_d : _GEN_279; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_474 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_d : _GEN_280; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_475 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_d : _GEN_281; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_476 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_d : _GEN_282; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_477 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_d : _GEN_283; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_494 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_g : _GEN_300; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_495 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_g : _GEN_301; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_496 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_g : _GEN_302; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_497 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_g : _GEN_303; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_498 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_g : _GEN_304; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_499 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_g : _GEN_305; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_500 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_g : _GEN_306; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_501 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_g : _GEN_307; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_502 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_g : _GEN_308; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_503 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_g : _GEN_309; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_504 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_g : _GEN_310; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_505 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_g : _GEN_311; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_506 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_g : _GEN_312; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_507 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_g : _GEN_313; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_508 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_g : _GEN_314; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_509 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_g : _GEN_315; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_510 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_u : _GEN_316; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_511 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_u : _GEN_317; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_512 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_u : _GEN_318; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_513 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_u : _GEN_319; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_514 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_u : _GEN_320; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_515 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_u : _GEN_321; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_516 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_u : _GEN_322; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_517 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_u : _GEN_323; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_518 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_u : _GEN_324; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_519 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_u : _GEN_325; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_520 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_u : _GEN_326; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_521 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_u : _GEN_327; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_522 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_u : _GEN_328; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_523 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_u : _GEN_329; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_524 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_u : _GEN_330; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_525 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_u : _GEN_331; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_526 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_x : _GEN_332; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_527 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_x : _GEN_333; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_528 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_x : _GEN_334; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_529 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_x : _GEN_335; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_530 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_x : _GEN_336; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_531 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_x : _GEN_337; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_532 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_x : _GEN_338; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_533 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_x : _GEN_339; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_534 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_x : _GEN_340; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_535 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_x : _GEN_341; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_536 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_x : _GEN_342; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_537 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_x : _GEN_343; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_538 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_x : _GEN_344; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_539 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_x : _GEN_345; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_540 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_x : _GEN_346; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_541 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_x : _GEN_347; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_542 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_w : _GEN_348; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_543 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_w : _GEN_349; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_544 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_w : _GEN_350; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_545 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_w : _GEN_351; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_546 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_w : _GEN_352; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_547 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_w : _GEN_353; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_548 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_w : _GEN_354; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_549 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_w : _GEN_355; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_550 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_w : _GEN_356; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_551 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_w : _GEN_357; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_552 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_w : _GEN_358; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_553 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_w : _GEN_359; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_554 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_w : _GEN_360; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_555 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_w : _GEN_361; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_556 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_w : _GEN_362; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_557 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_w : _GEN_363; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_558 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_r : _GEN_364; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_559 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_r : _GEN_365; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_560 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_r : _GEN_366; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_561 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_r : _GEN_367; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_562 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_r : _GEN_368; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_563 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_r : _GEN_369; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_564 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_r : _GEN_370; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_565 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_r : _GEN_371; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_566 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_r : _GEN_372; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_567 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_r : _GEN_373; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_568 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_r : _GEN_374; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_569 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_r : _GEN_375; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_570 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_r : _GEN_376; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_571 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_r : _GEN_377; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_572 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_r : _GEN_378; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_573 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_r : _GEN_379; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_574 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_flag_v : _GEN_380; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_575 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_flag_v : _GEN_381; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_576 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_flag_v : _GEN_382; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_577 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_flag_v : _GEN_383; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_578 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_flag_v : _GEN_384; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_579 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_flag_v : _GEN_385; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_580 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_flag_v : _GEN_386; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_581 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_flag_v : _GEN_387; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_582 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_flag_v : _GEN_388; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_583 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_flag_v : _GEN_389; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_584 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_flag_v : _GEN_390; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_585 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_flag_v : _GEN_391; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_586 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_flag_v : _GEN_392; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_587 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_flag_v : _GEN_393; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_588 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_flag_v : _GEN_394; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire  _GEN_589 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_flag_v : _GEN_395; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_590 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_ppn : _GEN_396; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_591 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_ppn : _GEN_397; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_592 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_ppn : _GEN_398; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_593 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_ppn : _GEN_399; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_594 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_ppn : _GEN_400; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_595 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_ppn : _GEN_401; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_596 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_ppn : _GEN_402; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_597 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_ppn : _GEN_403; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_598 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_ppn : _GEN_404; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_599 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_ppn : _GEN_405; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_600 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_ppn : _GEN_406; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_601 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_ppn : _GEN_407; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_602 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_ppn : _GEN_408; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_603 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_ppn : _GEN_409; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_604 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_ppn : _GEN_410; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [19:0] _GEN_605 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_ppn : _GEN_411; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_606 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_0_rmask : _GEN_412; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_607 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_1_rmask : _GEN_413; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_608 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_2_rmask : _GEN_414; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_609 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_3_rmask : _GEN_415; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_610 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_4_rmask : _GEN_416; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_611 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_5_rmask : _GEN_417; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_612 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_6_rmask : _GEN_418; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_613 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_7_rmask : _GEN_419; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_614 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_8_rmask : _GEN_420; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_615 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_9_rmask : _GEN_421; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_616 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_10_rmask : _GEN_422; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_617 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_11_rmask : _GEN_423; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_618 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_12_rmask : _GEN_424; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_619 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_13_rmask : _GEN_425; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_620 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_14_rmask : _GEN_426; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [17:0] _GEN_621 = io_dcache_ptw_pte_bits_page_fault ? tlbl2_15_rmask : _GEN_427; // @[playground/src/cache/mmu/Tlb.scala 236:55 77:22]
  wire [26:0] _GEN_622 = io_dcache_ptw_pte_bits_page_fault ? itlb_vpn : ivpn; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire [15:0] _GEN_623 = io_dcache_ptw_pte_bits_page_fault ? itlb_asid : satp_asid; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire  _GEN_626 = io_dcache_ptw_pte_bits_page_fault ? itlb_flag_g : io_dcache_ptw_pte_bits_entry_flag_g; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire  _GEN_627 = io_dcache_ptw_pte_bits_page_fault ? itlb_flag_u : io_dcache_ptw_pte_bits_entry_flag_u; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire  _GEN_628 = io_dcache_ptw_pte_bits_page_fault ? itlb_flag_x : io_dcache_ptw_pte_bits_entry_flag_x; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire  _GEN_631 = io_dcache_ptw_pte_bits_page_fault ? itlb_flag_v : io_dcache_ptw_pte_bits_entry_flag_v; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire [19:0] _GEN_632 = io_dcache_ptw_pte_bits_page_fault ? itlb_ppn : io_dcache_ptw_pte_bits_entry_ppn; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire [17:0] _GEN_633 = io_dcache_ptw_pte_bits_page_fault ? itlb_rmask : io_dcache_ptw_pte_bits_rmask; // @[playground/src/cache/mmu/Tlb.scala 236:55 75:22 248:38]
  wire [3:0] _GEN_634 = io_dcache_ptw_pte_bits_page_fault ? replace_index_value : _value_T_1; // @[playground/src/cache/mmu/Tlb.scala 236:55 src/main/scala/chisel3/util/Counter.scala 61:40 77:15]
  wire [1:0] _GEN_844 = io_dcache_ptw_pte_valid ? _GEN_429 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 232:37 106:76]
  wire  _GEN_845 = io_dcache_ptw_pte_valid ? _GEN_428 : ipage_fault; // @[playground/src/cache/mmu/Tlb.scala 112:30 232:37]
  wire [26:0] _GEN_846 = io_dcache_ptw_pte_valid ? _GEN_430 : tlbl2_0_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_847 = io_dcache_ptw_pte_valid ? _GEN_431 : tlbl2_1_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_848 = io_dcache_ptw_pte_valid ? _GEN_432 : tlbl2_2_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_849 = io_dcache_ptw_pte_valid ? _GEN_433 : tlbl2_3_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_850 = io_dcache_ptw_pte_valid ? _GEN_434 : tlbl2_4_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_851 = io_dcache_ptw_pte_valid ? _GEN_435 : tlbl2_5_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_852 = io_dcache_ptw_pte_valid ? _GEN_436 : tlbl2_6_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_853 = io_dcache_ptw_pte_valid ? _GEN_437 : tlbl2_7_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_854 = io_dcache_ptw_pte_valid ? _GEN_438 : tlbl2_8_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_855 = io_dcache_ptw_pte_valid ? _GEN_439 : tlbl2_9_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_856 = io_dcache_ptw_pte_valid ? _GEN_440 : tlbl2_10_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_857 = io_dcache_ptw_pte_valid ? _GEN_441 : tlbl2_11_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_858 = io_dcache_ptw_pte_valid ? _GEN_442 : tlbl2_12_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_859 = io_dcache_ptw_pte_valid ? _GEN_443 : tlbl2_13_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_860 = io_dcache_ptw_pte_valid ? _GEN_444 : tlbl2_14_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_861 = io_dcache_ptw_pte_valid ? _GEN_445 : tlbl2_15_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_862 = io_dcache_ptw_pte_valid ? _GEN_446 : tlbl2_0_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_863 = io_dcache_ptw_pte_valid ? _GEN_447 : tlbl2_1_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_864 = io_dcache_ptw_pte_valid ? _GEN_448 : tlbl2_2_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_865 = io_dcache_ptw_pte_valid ? _GEN_449 : tlbl2_3_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_866 = io_dcache_ptw_pte_valid ? _GEN_450 : tlbl2_4_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_867 = io_dcache_ptw_pte_valid ? _GEN_451 : tlbl2_5_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_868 = io_dcache_ptw_pte_valid ? _GEN_452 : tlbl2_6_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_869 = io_dcache_ptw_pte_valid ? _GEN_453 : tlbl2_7_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_870 = io_dcache_ptw_pte_valid ? _GEN_454 : tlbl2_8_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_871 = io_dcache_ptw_pte_valid ? _GEN_455 : tlbl2_9_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_872 = io_dcache_ptw_pte_valid ? _GEN_456 : tlbl2_10_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_873 = io_dcache_ptw_pte_valid ? _GEN_457 : tlbl2_11_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_874 = io_dcache_ptw_pte_valid ? _GEN_458 : tlbl2_12_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_875 = io_dcache_ptw_pte_valid ? _GEN_459 : tlbl2_13_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_876 = io_dcache_ptw_pte_valid ? _GEN_460 : tlbl2_14_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [15:0] _GEN_877 = io_dcache_ptw_pte_valid ? _GEN_461 : tlbl2_15_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_878 = io_dcache_ptw_pte_valid ? _GEN_462 : tlbl2_0_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_879 = io_dcache_ptw_pte_valid ? _GEN_463 : tlbl2_1_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_880 = io_dcache_ptw_pte_valid ? _GEN_464 : tlbl2_2_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_881 = io_dcache_ptw_pte_valid ? _GEN_465 : tlbl2_3_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_882 = io_dcache_ptw_pte_valid ? _GEN_466 : tlbl2_4_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_883 = io_dcache_ptw_pte_valid ? _GEN_467 : tlbl2_5_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_884 = io_dcache_ptw_pte_valid ? _GEN_468 : tlbl2_6_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_885 = io_dcache_ptw_pte_valid ? _GEN_469 : tlbl2_7_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_886 = io_dcache_ptw_pte_valid ? _GEN_470 : tlbl2_8_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_887 = io_dcache_ptw_pte_valid ? _GEN_471 : tlbl2_9_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_888 = io_dcache_ptw_pte_valid ? _GEN_472 : tlbl2_10_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_889 = io_dcache_ptw_pte_valid ? _GEN_473 : tlbl2_11_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_890 = io_dcache_ptw_pte_valid ? _GEN_474 : tlbl2_12_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_891 = io_dcache_ptw_pte_valid ? _GEN_475 : tlbl2_13_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_892 = io_dcache_ptw_pte_valid ? _GEN_476 : tlbl2_14_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_893 = io_dcache_ptw_pte_valid ? _GEN_477 : tlbl2_15_flag_d; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_910 = io_dcache_ptw_pte_valid ? _GEN_494 : tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_911 = io_dcache_ptw_pte_valid ? _GEN_495 : tlbl2_1_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_912 = io_dcache_ptw_pte_valid ? _GEN_496 : tlbl2_2_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_913 = io_dcache_ptw_pte_valid ? _GEN_497 : tlbl2_3_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_914 = io_dcache_ptw_pte_valid ? _GEN_498 : tlbl2_4_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_915 = io_dcache_ptw_pte_valid ? _GEN_499 : tlbl2_5_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_916 = io_dcache_ptw_pte_valid ? _GEN_500 : tlbl2_6_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_917 = io_dcache_ptw_pte_valid ? _GEN_501 : tlbl2_7_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_918 = io_dcache_ptw_pte_valid ? _GEN_502 : tlbl2_8_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_919 = io_dcache_ptw_pte_valid ? _GEN_503 : tlbl2_9_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_920 = io_dcache_ptw_pte_valid ? _GEN_504 : tlbl2_10_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_921 = io_dcache_ptw_pte_valid ? _GEN_505 : tlbl2_11_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_922 = io_dcache_ptw_pte_valid ? _GEN_506 : tlbl2_12_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_923 = io_dcache_ptw_pte_valid ? _GEN_507 : tlbl2_13_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_924 = io_dcache_ptw_pte_valid ? _GEN_508 : tlbl2_14_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_925 = io_dcache_ptw_pte_valid ? _GEN_509 : tlbl2_15_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_926 = io_dcache_ptw_pte_valid ? _GEN_510 : tlbl2_0_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_927 = io_dcache_ptw_pte_valid ? _GEN_511 : tlbl2_1_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_928 = io_dcache_ptw_pte_valid ? _GEN_512 : tlbl2_2_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_929 = io_dcache_ptw_pte_valid ? _GEN_513 : tlbl2_3_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_930 = io_dcache_ptw_pte_valid ? _GEN_514 : tlbl2_4_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_931 = io_dcache_ptw_pte_valid ? _GEN_515 : tlbl2_5_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_932 = io_dcache_ptw_pte_valid ? _GEN_516 : tlbl2_6_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_933 = io_dcache_ptw_pte_valid ? _GEN_517 : tlbl2_7_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_934 = io_dcache_ptw_pte_valid ? _GEN_518 : tlbl2_8_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_935 = io_dcache_ptw_pte_valid ? _GEN_519 : tlbl2_9_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_936 = io_dcache_ptw_pte_valid ? _GEN_520 : tlbl2_10_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_937 = io_dcache_ptw_pte_valid ? _GEN_521 : tlbl2_11_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_938 = io_dcache_ptw_pte_valid ? _GEN_522 : tlbl2_12_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_939 = io_dcache_ptw_pte_valid ? _GEN_523 : tlbl2_13_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_940 = io_dcache_ptw_pte_valid ? _GEN_524 : tlbl2_14_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_941 = io_dcache_ptw_pte_valid ? _GEN_525 : tlbl2_15_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_942 = io_dcache_ptw_pte_valid ? _GEN_526 : tlbl2_0_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_943 = io_dcache_ptw_pte_valid ? _GEN_527 : tlbl2_1_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_944 = io_dcache_ptw_pte_valid ? _GEN_528 : tlbl2_2_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_945 = io_dcache_ptw_pte_valid ? _GEN_529 : tlbl2_3_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_946 = io_dcache_ptw_pte_valid ? _GEN_530 : tlbl2_4_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_947 = io_dcache_ptw_pte_valid ? _GEN_531 : tlbl2_5_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_948 = io_dcache_ptw_pte_valid ? _GEN_532 : tlbl2_6_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_949 = io_dcache_ptw_pte_valid ? _GEN_533 : tlbl2_7_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_950 = io_dcache_ptw_pte_valid ? _GEN_534 : tlbl2_8_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_951 = io_dcache_ptw_pte_valid ? _GEN_535 : tlbl2_9_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_952 = io_dcache_ptw_pte_valid ? _GEN_536 : tlbl2_10_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_953 = io_dcache_ptw_pte_valid ? _GEN_537 : tlbl2_11_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_954 = io_dcache_ptw_pte_valid ? _GEN_538 : tlbl2_12_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_955 = io_dcache_ptw_pte_valid ? _GEN_539 : tlbl2_13_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_956 = io_dcache_ptw_pte_valid ? _GEN_540 : tlbl2_14_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_957 = io_dcache_ptw_pte_valid ? _GEN_541 : tlbl2_15_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_958 = io_dcache_ptw_pte_valid ? _GEN_542 : tlbl2_0_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_959 = io_dcache_ptw_pte_valid ? _GEN_543 : tlbl2_1_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_960 = io_dcache_ptw_pte_valid ? _GEN_544 : tlbl2_2_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_961 = io_dcache_ptw_pte_valid ? _GEN_545 : tlbl2_3_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_962 = io_dcache_ptw_pte_valid ? _GEN_546 : tlbl2_4_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_963 = io_dcache_ptw_pte_valid ? _GEN_547 : tlbl2_5_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_964 = io_dcache_ptw_pte_valid ? _GEN_548 : tlbl2_6_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_965 = io_dcache_ptw_pte_valid ? _GEN_549 : tlbl2_7_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_966 = io_dcache_ptw_pte_valid ? _GEN_550 : tlbl2_8_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_967 = io_dcache_ptw_pte_valid ? _GEN_551 : tlbl2_9_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_968 = io_dcache_ptw_pte_valid ? _GEN_552 : tlbl2_10_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_969 = io_dcache_ptw_pte_valid ? _GEN_553 : tlbl2_11_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_970 = io_dcache_ptw_pte_valid ? _GEN_554 : tlbl2_12_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_971 = io_dcache_ptw_pte_valid ? _GEN_555 : tlbl2_13_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_972 = io_dcache_ptw_pte_valid ? _GEN_556 : tlbl2_14_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_973 = io_dcache_ptw_pte_valid ? _GEN_557 : tlbl2_15_flag_w; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_974 = io_dcache_ptw_pte_valid ? _GEN_558 : tlbl2_0_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_975 = io_dcache_ptw_pte_valid ? _GEN_559 : tlbl2_1_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_976 = io_dcache_ptw_pte_valid ? _GEN_560 : tlbl2_2_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_977 = io_dcache_ptw_pte_valid ? _GEN_561 : tlbl2_3_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_978 = io_dcache_ptw_pte_valid ? _GEN_562 : tlbl2_4_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_979 = io_dcache_ptw_pte_valid ? _GEN_563 : tlbl2_5_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_980 = io_dcache_ptw_pte_valid ? _GEN_564 : tlbl2_6_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_981 = io_dcache_ptw_pte_valid ? _GEN_565 : tlbl2_7_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_982 = io_dcache_ptw_pte_valid ? _GEN_566 : tlbl2_8_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_983 = io_dcache_ptw_pte_valid ? _GEN_567 : tlbl2_9_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_984 = io_dcache_ptw_pte_valid ? _GEN_568 : tlbl2_10_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_985 = io_dcache_ptw_pte_valid ? _GEN_569 : tlbl2_11_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_986 = io_dcache_ptw_pte_valid ? _GEN_570 : tlbl2_12_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_987 = io_dcache_ptw_pte_valid ? _GEN_571 : tlbl2_13_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_988 = io_dcache_ptw_pte_valid ? _GEN_572 : tlbl2_14_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_989 = io_dcache_ptw_pte_valid ? _GEN_573 : tlbl2_15_flag_r; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_990 = io_dcache_ptw_pte_valid ? _GEN_574 : tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_991 = io_dcache_ptw_pte_valid ? _GEN_575 : tlbl2_1_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_992 = io_dcache_ptw_pte_valid ? _GEN_576 : tlbl2_2_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_993 = io_dcache_ptw_pte_valid ? _GEN_577 : tlbl2_3_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_994 = io_dcache_ptw_pte_valid ? _GEN_578 : tlbl2_4_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_995 = io_dcache_ptw_pte_valid ? _GEN_579 : tlbl2_5_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_996 = io_dcache_ptw_pte_valid ? _GEN_580 : tlbl2_6_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_997 = io_dcache_ptw_pte_valid ? _GEN_581 : tlbl2_7_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_998 = io_dcache_ptw_pte_valid ? _GEN_582 : tlbl2_8_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_999 = io_dcache_ptw_pte_valid ? _GEN_583 : tlbl2_9_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_1000 = io_dcache_ptw_pte_valid ? _GEN_584 : tlbl2_10_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_1001 = io_dcache_ptw_pte_valid ? _GEN_585 : tlbl2_11_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_1002 = io_dcache_ptw_pte_valid ? _GEN_586 : tlbl2_12_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_1003 = io_dcache_ptw_pte_valid ? _GEN_587 : tlbl2_13_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_1004 = io_dcache_ptw_pte_valid ? _GEN_588 : tlbl2_14_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire  _GEN_1005 = io_dcache_ptw_pte_valid ? _GEN_589 : tlbl2_15_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1006 = io_dcache_ptw_pte_valid ? _GEN_590 : tlbl2_0_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1007 = io_dcache_ptw_pte_valid ? _GEN_591 : tlbl2_1_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1008 = io_dcache_ptw_pte_valid ? _GEN_592 : tlbl2_2_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1009 = io_dcache_ptw_pte_valid ? _GEN_593 : tlbl2_3_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1010 = io_dcache_ptw_pte_valid ? _GEN_594 : tlbl2_4_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1011 = io_dcache_ptw_pte_valid ? _GEN_595 : tlbl2_5_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1012 = io_dcache_ptw_pte_valid ? _GEN_596 : tlbl2_6_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1013 = io_dcache_ptw_pte_valid ? _GEN_597 : tlbl2_7_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1014 = io_dcache_ptw_pte_valid ? _GEN_598 : tlbl2_8_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1015 = io_dcache_ptw_pte_valid ? _GEN_599 : tlbl2_9_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1016 = io_dcache_ptw_pte_valid ? _GEN_600 : tlbl2_10_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1017 = io_dcache_ptw_pte_valid ? _GEN_601 : tlbl2_11_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1018 = io_dcache_ptw_pte_valid ? _GEN_602 : tlbl2_12_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1019 = io_dcache_ptw_pte_valid ? _GEN_603 : tlbl2_13_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1020 = io_dcache_ptw_pte_valid ? _GEN_604 : tlbl2_14_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [19:0] _GEN_1021 = io_dcache_ptw_pte_valid ? _GEN_605 : tlbl2_15_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1022 = io_dcache_ptw_pte_valid ? _GEN_606 : tlbl2_0_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1023 = io_dcache_ptw_pte_valid ? _GEN_607 : tlbl2_1_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1024 = io_dcache_ptw_pte_valid ? _GEN_608 : tlbl2_2_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1025 = io_dcache_ptw_pte_valid ? _GEN_609 : tlbl2_3_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1026 = io_dcache_ptw_pte_valid ? _GEN_610 : tlbl2_4_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1027 = io_dcache_ptw_pte_valid ? _GEN_611 : tlbl2_5_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1028 = io_dcache_ptw_pte_valid ? _GEN_612 : tlbl2_6_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1029 = io_dcache_ptw_pte_valid ? _GEN_613 : tlbl2_7_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1030 = io_dcache_ptw_pte_valid ? _GEN_614 : tlbl2_8_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1031 = io_dcache_ptw_pte_valid ? _GEN_615 : tlbl2_9_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1032 = io_dcache_ptw_pte_valid ? _GEN_616 : tlbl2_10_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1033 = io_dcache_ptw_pte_valid ? _GEN_617 : tlbl2_11_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1034 = io_dcache_ptw_pte_valid ? _GEN_618 : tlbl2_12_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1035 = io_dcache_ptw_pte_valid ? _GEN_619 : tlbl2_13_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1036 = io_dcache_ptw_pte_valid ? _GEN_620 : tlbl2_14_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [17:0] _GEN_1037 = io_dcache_ptw_pte_valid ? _GEN_621 : tlbl2_15_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 77:22]
  wire [26:0] _GEN_1038 = io_dcache_ptw_pte_valid ? _GEN_622 : itlb_vpn; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire [15:0] _GEN_1039 = io_dcache_ptw_pte_valid ? _GEN_623 : itlb_asid; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire  _GEN_1042 = io_dcache_ptw_pte_valid ? _GEN_626 : itlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire  _GEN_1043 = io_dcache_ptw_pte_valid ? _GEN_627 : itlb_flag_u; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire  _GEN_1044 = io_dcache_ptw_pte_valid ? _GEN_628 : itlb_flag_x; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire  _GEN_1047 = io_dcache_ptw_pte_valid ? _GEN_631 : itlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire [19:0] _GEN_1048 = io_dcache_ptw_pte_valid ? _GEN_632 : itlb_ppn; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire [17:0] _GEN_1049 = io_dcache_ptw_pte_valid ? _GEN_633 : itlb_rmask; // @[playground/src/cache/mmu/Tlb.scala 232:37 75:22]
  wire [3:0] _GEN_1050 = io_dcache_ptw_pte_valid ? _GEN_634 : replace_index_value; // @[playground/src/cache/mmu/Tlb.scala 232:37 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _GEN_1051 = io_icache_complete_single_request ? 1'h0 : ipage_fault; // @[playground/src/cache/mmu/Tlb.scala 255:47 256:23 112:30]
  wire [1:0] _GEN_1053 = io_icache_complete_single_request ? 2'h0 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 255:47 258:23 106:76]
  wire  _GEN_1054 = 2'h3 == immu_state ? _GEN_1051 : ipage_fault; // @[playground/src/cache/mmu/Tlb.scala 193:22 112:30]
  wire [1:0] _GEN_1056 = 2'h3 == immu_state ? _GEN_1053 : immu_state; // @[playground/src/cache/mmu/Tlb.scala 193:22 106:76]
  wire [26:0] _GEN_1061 = 2'h2 == immu_state ? _GEN_846 : tlbl2_0_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1062 = 2'h2 == immu_state ? _GEN_847 : tlbl2_1_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1063 = 2'h2 == immu_state ? _GEN_848 : tlbl2_2_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1064 = 2'h2 == immu_state ? _GEN_849 : tlbl2_3_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1065 = 2'h2 == immu_state ? _GEN_850 : tlbl2_4_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1066 = 2'h2 == immu_state ? _GEN_851 : tlbl2_5_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1067 = 2'h2 == immu_state ? _GEN_852 : tlbl2_6_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1068 = 2'h2 == immu_state ? _GEN_853 : tlbl2_7_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1069 = 2'h2 == immu_state ? _GEN_854 : tlbl2_8_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1070 = 2'h2 == immu_state ? _GEN_855 : tlbl2_9_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1071 = 2'h2 == immu_state ? _GEN_856 : tlbl2_10_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1072 = 2'h2 == immu_state ? _GEN_857 : tlbl2_11_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1073 = 2'h2 == immu_state ? _GEN_858 : tlbl2_12_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1074 = 2'h2 == immu_state ? _GEN_859 : tlbl2_13_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1075 = 2'h2 == immu_state ? _GEN_860 : tlbl2_14_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1076 = 2'h2 == immu_state ? _GEN_861 : tlbl2_15_vpn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1077 = 2'h2 == immu_state ? _GEN_862 : tlbl2_0_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1078 = 2'h2 == immu_state ? _GEN_863 : tlbl2_1_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1079 = 2'h2 == immu_state ? _GEN_864 : tlbl2_2_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1080 = 2'h2 == immu_state ? _GEN_865 : tlbl2_3_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1081 = 2'h2 == immu_state ? _GEN_866 : tlbl2_4_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1082 = 2'h2 == immu_state ? _GEN_867 : tlbl2_5_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1083 = 2'h2 == immu_state ? _GEN_868 : tlbl2_6_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1084 = 2'h2 == immu_state ? _GEN_869 : tlbl2_7_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1085 = 2'h2 == immu_state ? _GEN_870 : tlbl2_8_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1086 = 2'h2 == immu_state ? _GEN_871 : tlbl2_9_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1087 = 2'h2 == immu_state ? _GEN_872 : tlbl2_10_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1088 = 2'h2 == immu_state ? _GEN_873 : tlbl2_11_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1089 = 2'h2 == immu_state ? _GEN_874 : tlbl2_12_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1090 = 2'h2 == immu_state ? _GEN_875 : tlbl2_13_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1091 = 2'h2 == immu_state ? _GEN_876 : tlbl2_14_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1092 = 2'h2 == immu_state ? _GEN_877 : tlbl2_15_asid; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1093 = 2'h2 == immu_state ? _GEN_878 : tlbl2_0_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1094 = 2'h2 == immu_state ? _GEN_879 : tlbl2_1_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1095 = 2'h2 == immu_state ? _GEN_880 : tlbl2_2_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1096 = 2'h2 == immu_state ? _GEN_881 : tlbl2_3_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1097 = 2'h2 == immu_state ? _GEN_882 : tlbl2_4_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1098 = 2'h2 == immu_state ? _GEN_883 : tlbl2_5_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1099 = 2'h2 == immu_state ? _GEN_884 : tlbl2_6_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1100 = 2'h2 == immu_state ? _GEN_885 : tlbl2_7_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1101 = 2'h2 == immu_state ? _GEN_886 : tlbl2_8_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1102 = 2'h2 == immu_state ? _GEN_887 : tlbl2_9_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1103 = 2'h2 == immu_state ? _GEN_888 : tlbl2_10_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1104 = 2'h2 == immu_state ? _GEN_889 : tlbl2_11_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1105 = 2'h2 == immu_state ? _GEN_890 : tlbl2_12_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1106 = 2'h2 == immu_state ? _GEN_891 : tlbl2_13_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1107 = 2'h2 == immu_state ? _GEN_892 : tlbl2_14_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1108 = 2'h2 == immu_state ? _GEN_893 : tlbl2_15_flag_d; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1125 = 2'h2 == immu_state ? _GEN_910 : tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1126 = 2'h2 == immu_state ? _GEN_911 : tlbl2_1_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1127 = 2'h2 == immu_state ? _GEN_912 : tlbl2_2_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1128 = 2'h2 == immu_state ? _GEN_913 : tlbl2_3_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1129 = 2'h2 == immu_state ? _GEN_914 : tlbl2_4_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1130 = 2'h2 == immu_state ? _GEN_915 : tlbl2_5_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1131 = 2'h2 == immu_state ? _GEN_916 : tlbl2_6_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1132 = 2'h2 == immu_state ? _GEN_917 : tlbl2_7_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1133 = 2'h2 == immu_state ? _GEN_918 : tlbl2_8_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1134 = 2'h2 == immu_state ? _GEN_919 : tlbl2_9_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1135 = 2'h2 == immu_state ? _GEN_920 : tlbl2_10_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1136 = 2'h2 == immu_state ? _GEN_921 : tlbl2_11_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1137 = 2'h2 == immu_state ? _GEN_922 : tlbl2_12_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1138 = 2'h2 == immu_state ? _GEN_923 : tlbl2_13_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1139 = 2'h2 == immu_state ? _GEN_924 : tlbl2_14_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1140 = 2'h2 == immu_state ? _GEN_925 : tlbl2_15_flag_g; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1141 = 2'h2 == immu_state ? _GEN_926 : tlbl2_0_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1142 = 2'h2 == immu_state ? _GEN_927 : tlbl2_1_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1143 = 2'h2 == immu_state ? _GEN_928 : tlbl2_2_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1144 = 2'h2 == immu_state ? _GEN_929 : tlbl2_3_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1145 = 2'h2 == immu_state ? _GEN_930 : tlbl2_4_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1146 = 2'h2 == immu_state ? _GEN_931 : tlbl2_5_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1147 = 2'h2 == immu_state ? _GEN_932 : tlbl2_6_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1148 = 2'h2 == immu_state ? _GEN_933 : tlbl2_7_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1149 = 2'h2 == immu_state ? _GEN_934 : tlbl2_8_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1150 = 2'h2 == immu_state ? _GEN_935 : tlbl2_9_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1151 = 2'h2 == immu_state ? _GEN_936 : tlbl2_10_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1152 = 2'h2 == immu_state ? _GEN_937 : tlbl2_11_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1153 = 2'h2 == immu_state ? _GEN_938 : tlbl2_12_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1154 = 2'h2 == immu_state ? _GEN_939 : tlbl2_13_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1155 = 2'h2 == immu_state ? _GEN_940 : tlbl2_14_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1156 = 2'h2 == immu_state ? _GEN_941 : tlbl2_15_flag_u; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1157 = 2'h2 == immu_state ? _GEN_942 : tlbl2_0_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1158 = 2'h2 == immu_state ? _GEN_943 : tlbl2_1_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1159 = 2'h2 == immu_state ? _GEN_944 : tlbl2_2_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1160 = 2'h2 == immu_state ? _GEN_945 : tlbl2_3_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1161 = 2'h2 == immu_state ? _GEN_946 : tlbl2_4_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1162 = 2'h2 == immu_state ? _GEN_947 : tlbl2_5_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1163 = 2'h2 == immu_state ? _GEN_948 : tlbl2_6_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1164 = 2'h2 == immu_state ? _GEN_949 : tlbl2_7_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1165 = 2'h2 == immu_state ? _GEN_950 : tlbl2_8_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1166 = 2'h2 == immu_state ? _GEN_951 : tlbl2_9_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1167 = 2'h2 == immu_state ? _GEN_952 : tlbl2_10_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1168 = 2'h2 == immu_state ? _GEN_953 : tlbl2_11_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1169 = 2'h2 == immu_state ? _GEN_954 : tlbl2_12_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1170 = 2'h2 == immu_state ? _GEN_955 : tlbl2_13_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1171 = 2'h2 == immu_state ? _GEN_956 : tlbl2_14_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1172 = 2'h2 == immu_state ? _GEN_957 : tlbl2_15_flag_x; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1173 = 2'h2 == immu_state ? _GEN_958 : tlbl2_0_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1174 = 2'h2 == immu_state ? _GEN_959 : tlbl2_1_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1175 = 2'h2 == immu_state ? _GEN_960 : tlbl2_2_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1176 = 2'h2 == immu_state ? _GEN_961 : tlbl2_3_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1177 = 2'h2 == immu_state ? _GEN_962 : tlbl2_4_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1178 = 2'h2 == immu_state ? _GEN_963 : tlbl2_5_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1179 = 2'h2 == immu_state ? _GEN_964 : tlbl2_6_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1180 = 2'h2 == immu_state ? _GEN_965 : tlbl2_7_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1181 = 2'h2 == immu_state ? _GEN_966 : tlbl2_8_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1182 = 2'h2 == immu_state ? _GEN_967 : tlbl2_9_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1183 = 2'h2 == immu_state ? _GEN_968 : tlbl2_10_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1184 = 2'h2 == immu_state ? _GEN_969 : tlbl2_11_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1185 = 2'h2 == immu_state ? _GEN_970 : tlbl2_12_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1186 = 2'h2 == immu_state ? _GEN_971 : tlbl2_13_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1187 = 2'h2 == immu_state ? _GEN_972 : tlbl2_14_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1188 = 2'h2 == immu_state ? _GEN_973 : tlbl2_15_flag_w; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1189 = 2'h2 == immu_state ? _GEN_974 : tlbl2_0_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1190 = 2'h2 == immu_state ? _GEN_975 : tlbl2_1_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1191 = 2'h2 == immu_state ? _GEN_976 : tlbl2_2_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1192 = 2'h2 == immu_state ? _GEN_977 : tlbl2_3_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1193 = 2'h2 == immu_state ? _GEN_978 : tlbl2_4_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1194 = 2'h2 == immu_state ? _GEN_979 : tlbl2_5_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1195 = 2'h2 == immu_state ? _GEN_980 : tlbl2_6_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1196 = 2'h2 == immu_state ? _GEN_981 : tlbl2_7_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1197 = 2'h2 == immu_state ? _GEN_982 : tlbl2_8_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1198 = 2'h2 == immu_state ? _GEN_983 : tlbl2_9_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1199 = 2'h2 == immu_state ? _GEN_984 : tlbl2_10_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1200 = 2'h2 == immu_state ? _GEN_985 : tlbl2_11_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1201 = 2'h2 == immu_state ? _GEN_986 : tlbl2_12_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1202 = 2'h2 == immu_state ? _GEN_987 : tlbl2_13_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1203 = 2'h2 == immu_state ? _GEN_988 : tlbl2_14_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1204 = 2'h2 == immu_state ? _GEN_989 : tlbl2_15_flag_r; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1205 = 2'h2 == immu_state ? _GEN_990 : tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1206 = 2'h2 == immu_state ? _GEN_991 : tlbl2_1_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1207 = 2'h2 == immu_state ? _GEN_992 : tlbl2_2_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1208 = 2'h2 == immu_state ? _GEN_993 : tlbl2_3_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1209 = 2'h2 == immu_state ? _GEN_994 : tlbl2_4_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1210 = 2'h2 == immu_state ? _GEN_995 : tlbl2_5_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1211 = 2'h2 == immu_state ? _GEN_996 : tlbl2_6_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1212 = 2'h2 == immu_state ? _GEN_997 : tlbl2_7_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1213 = 2'h2 == immu_state ? _GEN_998 : tlbl2_8_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1214 = 2'h2 == immu_state ? _GEN_999 : tlbl2_9_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1215 = 2'h2 == immu_state ? _GEN_1000 : tlbl2_10_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1216 = 2'h2 == immu_state ? _GEN_1001 : tlbl2_11_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1217 = 2'h2 == immu_state ? _GEN_1002 : tlbl2_12_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1218 = 2'h2 == immu_state ? _GEN_1003 : tlbl2_13_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1219 = 2'h2 == immu_state ? _GEN_1004 : tlbl2_14_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1220 = 2'h2 == immu_state ? _GEN_1005 : tlbl2_15_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1221 = 2'h2 == immu_state ? _GEN_1006 : tlbl2_0_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1222 = 2'h2 == immu_state ? _GEN_1007 : tlbl2_1_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1223 = 2'h2 == immu_state ? _GEN_1008 : tlbl2_2_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1224 = 2'h2 == immu_state ? _GEN_1009 : tlbl2_3_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1225 = 2'h2 == immu_state ? _GEN_1010 : tlbl2_4_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1226 = 2'h2 == immu_state ? _GEN_1011 : tlbl2_5_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1227 = 2'h2 == immu_state ? _GEN_1012 : tlbl2_6_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1228 = 2'h2 == immu_state ? _GEN_1013 : tlbl2_7_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1229 = 2'h2 == immu_state ? _GEN_1014 : tlbl2_8_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1230 = 2'h2 == immu_state ? _GEN_1015 : tlbl2_9_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1231 = 2'h2 == immu_state ? _GEN_1016 : tlbl2_10_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1232 = 2'h2 == immu_state ? _GEN_1017 : tlbl2_11_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1233 = 2'h2 == immu_state ? _GEN_1018 : tlbl2_12_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1234 = 2'h2 == immu_state ? _GEN_1019 : tlbl2_13_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1235 = 2'h2 == immu_state ? _GEN_1020 : tlbl2_14_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1236 = 2'h2 == immu_state ? _GEN_1021 : tlbl2_15_ppn; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1237 = 2'h2 == immu_state ? _GEN_1022 : tlbl2_0_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1238 = 2'h2 == immu_state ? _GEN_1023 : tlbl2_1_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1239 = 2'h2 == immu_state ? _GEN_1024 : tlbl2_2_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1240 = 2'h2 == immu_state ? _GEN_1025 : tlbl2_3_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1241 = 2'h2 == immu_state ? _GEN_1026 : tlbl2_4_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1242 = 2'h2 == immu_state ? _GEN_1027 : tlbl2_5_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1243 = 2'h2 == immu_state ? _GEN_1028 : tlbl2_6_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1244 = 2'h2 == immu_state ? _GEN_1029 : tlbl2_7_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1245 = 2'h2 == immu_state ? _GEN_1030 : tlbl2_8_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1246 = 2'h2 == immu_state ? _GEN_1031 : tlbl2_9_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1247 = 2'h2 == immu_state ? _GEN_1032 : tlbl2_10_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1248 = 2'h2 == immu_state ? _GEN_1033 : tlbl2_11_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1249 = 2'h2 == immu_state ? _GEN_1034 : tlbl2_12_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1250 = 2'h2 == immu_state ? _GEN_1035 : tlbl2_13_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1251 = 2'h2 == immu_state ? _GEN_1036 : tlbl2_14_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1252 = 2'h2 == immu_state ? _GEN_1037 : tlbl2_15_rmask; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1262 = 2'h2 == immu_state ? _GEN_1047 : itlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 193:22 75:22]
  wire [3:0] _GEN_1265 = 2'h2 == immu_state ? _GEN_1050 : replace_index_value; // @[playground/src/cache/mmu/Tlb.scala 193:22 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _GEN_1276 = 2'h1 == immu_state ? _GEN_232 : _GEN_1262; // @[playground/src/cache/mmu/Tlb.scala 193:22]
  wire [26:0] _GEN_1282 = 2'h1 == immu_state ? tlbl2_0_vpn : _GEN_1061; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1283 = 2'h1 == immu_state ? tlbl2_1_vpn : _GEN_1062; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1284 = 2'h1 == immu_state ? tlbl2_2_vpn : _GEN_1063; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1285 = 2'h1 == immu_state ? tlbl2_3_vpn : _GEN_1064; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1286 = 2'h1 == immu_state ? tlbl2_4_vpn : _GEN_1065; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1287 = 2'h1 == immu_state ? tlbl2_5_vpn : _GEN_1066; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1288 = 2'h1 == immu_state ? tlbl2_6_vpn : _GEN_1067; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1289 = 2'h1 == immu_state ? tlbl2_7_vpn : _GEN_1068; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1290 = 2'h1 == immu_state ? tlbl2_8_vpn : _GEN_1069; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1291 = 2'h1 == immu_state ? tlbl2_9_vpn : _GEN_1070; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1292 = 2'h1 == immu_state ? tlbl2_10_vpn : _GEN_1071; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1293 = 2'h1 == immu_state ? tlbl2_11_vpn : _GEN_1072; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1294 = 2'h1 == immu_state ? tlbl2_12_vpn : _GEN_1073; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1295 = 2'h1 == immu_state ? tlbl2_13_vpn : _GEN_1074; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1296 = 2'h1 == immu_state ? tlbl2_14_vpn : _GEN_1075; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1297 = 2'h1 == immu_state ? tlbl2_15_vpn : _GEN_1076; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1298 = 2'h1 == immu_state ? tlbl2_0_asid : _GEN_1077; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1299 = 2'h1 == immu_state ? tlbl2_1_asid : _GEN_1078; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1300 = 2'h1 == immu_state ? tlbl2_2_asid : _GEN_1079; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1301 = 2'h1 == immu_state ? tlbl2_3_asid : _GEN_1080; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1302 = 2'h1 == immu_state ? tlbl2_4_asid : _GEN_1081; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1303 = 2'h1 == immu_state ? tlbl2_5_asid : _GEN_1082; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1304 = 2'h1 == immu_state ? tlbl2_6_asid : _GEN_1083; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1305 = 2'h1 == immu_state ? tlbl2_7_asid : _GEN_1084; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1306 = 2'h1 == immu_state ? tlbl2_8_asid : _GEN_1085; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1307 = 2'h1 == immu_state ? tlbl2_9_asid : _GEN_1086; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1308 = 2'h1 == immu_state ? tlbl2_10_asid : _GEN_1087; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1309 = 2'h1 == immu_state ? tlbl2_11_asid : _GEN_1088; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1310 = 2'h1 == immu_state ? tlbl2_12_asid : _GEN_1089; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1311 = 2'h1 == immu_state ? tlbl2_13_asid : _GEN_1090; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1312 = 2'h1 == immu_state ? tlbl2_14_asid : _GEN_1091; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1313 = 2'h1 == immu_state ? tlbl2_15_asid : _GEN_1092; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1314 = 2'h1 == immu_state ? tlbl2_0_flag_d : _GEN_1093; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1315 = 2'h1 == immu_state ? tlbl2_1_flag_d : _GEN_1094; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1316 = 2'h1 == immu_state ? tlbl2_2_flag_d : _GEN_1095; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1317 = 2'h1 == immu_state ? tlbl2_3_flag_d : _GEN_1096; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1318 = 2'h1 == immu_state ? tlbl2_4_flag_d : _GEN_1097; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1319 = 2'h1 == immu_state ? tlbl2_5_flag_d : _GEN_1098; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1320 = 2'h1 == immu_state ? tlbl2_6_flag_d : _GEN_1099; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1321 = 2'h1 == immu_state ? tlbl2_7_flag_d : _GEN_1100; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1322 = 2'h1 == immu_state ? tlbl2_8_flag_d : _GEN_1101; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1323 = 2'h1 == immu_state ? tlbl2_9_flag_d : _GEN_1102; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1324 = 2'h1 == immu_state ? tlbl2_10_flag_d : _GEN_1103; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1325 = 2'h1 == immu_state ? tlbl2_11_flag_d : _GEN_1104; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1326 = 2'h1 == immu_state ? tlbl2_12_flag_d : _GEN_1105; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1327 = 2'h1 == immu_state ? tlbl2_13_flag_d : _GEN_1106; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1328 = 2'h1 == immu_state ? tlbl2_14_flag_d : _GEN_1107; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1329 = 2'h1 == immu_state ? tlbl2_15_flag_d : _GEN_1108; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1346 = 2'h1 == immu_state ? tlbl2_0_flag_g : _GEN_1125; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1347 = 2'h1 == immu_state ? tlbl2_1_flag_g : _GEN_1126; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1348 = 2'h1 == immu_state ? tlbl2_2_flag_g : _GEN_1127; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1349 = 2'h1 == immu_state ? tlbl2_3_flag_g : _GEN_1128; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1350 = 2'h1 == immu_state ? tlbl2_4_flag_g : _GEN_1129; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1351 = 2'h1 == immu_state ? tlbl2_5_flag_g : _GEN_1130; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1352 = 2'h1 == immu_state ? tlbl2_6_flag_g : _GEN_1131; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1353 = 2'h1 == immu_state ? tlbl2_7_flag_g : _GEN_1132; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1354 = 2'h1 == immu_state ? tlbl2_8_flag_g : _GEN_1133; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1355 = 2'h1 == immu_state ? tlbl2_9_flag_g : _GEN_1134; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1356 = 2'h1 == immu_state ? tlbl2_10_flag_g : _GEN_1135; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1357 = 2'h1 == immu_state ? tlbl2_11_flag_g : _GEN_1136; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1358 = 2'h1 == immu_state ? tlbl2_12_flag_g : _GEN_1137; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1359 = 2'h1 == immu_state ? tlbl2_13_flag_g : _GEN_1138; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1360 = 2'h1 == immu_state ? tlbl2_14_flag_g : _GEN_1139; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1361 = 2'h1 == immu_state ? tlbl2_15_flag_g : _GEN_1140; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1362 = 2'h1 == immu_state ? tlbl2_0_flag_u : _GEN_1141; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1363 = 2'h1 == immu_state ? tlbl2_1_flag_u : _GEN_1142; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1364 = 2'h1 == immu_state ? tlbl2_2_flag_u : _GEN_1143; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1365 = 2'h1 == immu_state ? tlbl2_3_flag_u : _GEN_1144; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1366 = 2'h1 == immu_state ? tlbl2_4_flag_u : _GEN_1145; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1367 = 2'h1 == immu_state ? tlbl2_5_flag_u : _GEN_1146; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1368 = 2'h1 == immu_state ? tlbl2_6_flag_u : _GEN_1147; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1369 = 2'h1 == immu_state ? tlbl2_7_flag_u : _GEN_1148; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1370 = 2'h1 == immu_state ? tlbl2_8_flag_u : _GEN_1149; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1371 = 2'h1 == immu_state ? tlbl2_9_flag_u : _GEN_1150; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1372 = 2'h1 == immu_state ? tlbl2_10_flag_u : _GEN_1151; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1373 = 2'h1 == immu_state ? tlbl2_11_flag_u : _GEN_1152; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1374 = 2'h1 == immu_state ? tlbl2_12_flag_u : _GEN_1153; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1375 = 2'h1 == immu_state ? tlbl2_13_flag_u : _GEN_1154; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1376 = 2'h1 == immu_state ? tlbl2_14_flag_u : _GEN_1155; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1377 = 2'h1 == immu_state ? tlbl2_15_flag_u : _GEN_1156; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1378 = 2'h1 == immu_state ? tlbl2_0_flag_x : _GEN_1157; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1379 = 2'h1 == immu_state ? tlbl2_1_flag_x : _GEN_1158; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1380 = 2'h1 == immu_state ? tlbl2_2_flag_x : _GEN_1159; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1381 = 2'h1 == immu_state ? tlbl2_3_flag_x : _GEN_1160; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1382 = 2'h1 == immu_state ? tlbl2_4_flag_x : _GEN_1161; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1383 = 2'h1 == immu_state ? tlbl2_5_flag_x : _GEN_1162; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1384 = 2'h1 == immu_state ? tlbl2_6_flag_x : _GEN_1163; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1385 = 2'h1 == immu_state ? tlbl2_7_flag_x : _GEN_1164; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1386 = 2'h1 == immu_state ? tlbl2_8_flag_x : _GEN_1165; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1387 = 2'h1 == immu_state ? tlbl2_9_flag_x : _GEN_1166; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1388 = 2'h1 == immu_state ? tlbl2_10_flag_x : _GEN_1167; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1389 = 2'h1 == immu_state ? tlbl2_11_flag_x : _GEN_1168; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1390 = 2'h1 == immu_state ? tlbl2_12_flag_x : _GEN_1169; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1391 = 2'h1 == immu_state ? tlbl2_13_flag_x : _GEN_1170; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1392 = 2'h1 == immu_state ? tlbl2_14_flag_x : _GEN_1171; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1393 = 2'h1 == immu_state ? tlbl2_15_flag_x : _GEN_1172; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1394 = 2'h1 == immu_state ? tlbl2_0_flag_w : _GEN_1173; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1395 = 2'h1 == immu_state ? tlbl2_1_flag_w : _GEN_1174; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1396 = 2'h1 == immu_state ? tlbl2_2_flag_w : _GEN_1175; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1397 = 2'h1 == immu_state ? tlbl2_3_flag_w : _GEN_1176; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1398 = 2'h1 == immu_state ? tlbl2_4_flag_w : _GEN_1177; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1399 = 2'h1 == immu_state ? tlbl2_5_flag_w : _GEN_1178; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1400 = 2'h1 == immu_state ? tlbl2_6_flag_w : _GEN_1179; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1401 = 2'h1 == immu_state ? tlbl2_7_flag_w : _GEN_1180; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1402 = 2'h1 == immu_state ? tlbl2_8_flag_w : _GEN_1181; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1403 = 2'h1 == immu_state ? tlbl2_9_flag_w : _GEN_1182; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1404 = 2'h1 == immu_state ? tlbl2_10_flag_w : _GEN_1183; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1405 = 2'h1 == immu_state ? tlbl2_11_flag_w : _GEN_1184; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1406 = 2'h1 == immu_state ? tlbl2_12_flag_w : _GEN_1185; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1407 = 2'h1 == immu_state ? tlbl2_13_flag_w : _GEN_1186; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1408 = 2'h1 == immu_state ? tlbl2_14_flag_w : _GEN_1187; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1409 = 2'h1 == immu_state ? tlbl2_15_flag_w : _GEN_1188; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1410 = 2'h1 == immu_state ? tlbl2_0_flag_r : _GEN_1189; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1411 = 2'h1 == immu_state ? tlbl2_1_flag_r : _GEN_1190; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1412 = 2'h1 == immu_state ? tlbl2_2_flag_r : _GEN_1191; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1413 = 2'h1 == immu_state ? tlbl2_3_flag_r : _GEN_1192; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1414 = 2'h1 == immu_state ? tlbl2_4_flag_r : _GEN_1193; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1415 = 2'h1 == immu_state ? tlbl2_5_flag_r : _GEN_1194; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1416 = 2'h1 == immu_state ? tlbl2_6_flag_r : _GEN_1195; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1417 = 2'h1 == immu_state ? tlbl2_7_flag_r : _GEN_1196; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1418 = 2'h1 == immu_state ? tlbl2_8_flag_r : _GEN_1197; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1419 = 2'h1 == immu_state ? tlbl2_9_flag_r : _GEN_1198; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1420 = 2'h1 == immu_state ? tlbl2_10_flag_r : _GEN_1199; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1421 = 2'h1 == immu_state ? tlbl2_11_flag_r : _GEN_1200; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1422 = 2'h1 == immu_state ? tlbl2_12_flag_r : _GEN_1201; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1423 = 2'h1 == immu_state ? tlbl2_13_flag_r : _GEN_1202; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1424 = 2'h1 == immu_state ? tlbl2_14_flag_r : _GEN_1203; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1425 = 2'h1 == immu_state ? tlbl2_15_flag_r : _GEN_1204; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1426 = 2'h1 == immu_state ? tlbl2_0_flag_v : _GEN_1205; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1427 = 2'h1 == immu_state ? tlbl2_1_flag_v : _GEN_1206; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1428 = 2'h1 == immu_state ? tlbl2_2_flag_v : _GEN_1207; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1429 = 2'h1 == immu_state ? tlbl2_3_flag_v : _GEN_1208; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1430 = 2'h1 == immu_state ? tlbl2_4_flag_v : _GEN_1209; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1431 = 2'h1 == immu_state ? tlbl2_5_flag_v : _GEN_1210; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1432 = 2'h1 == immu_state ? tlbl2_6_flag_v : _GEN_1211; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1433 = 2'h1 == immu_state ? tlbl2_7_flag_v : _GEN_1212; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1434 = 2'h1 == immu_state ? tlbl2_8_flag_v : _GEN_1213; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1435 = 2'h1 == immu_state ? tlbl2_9_flag_v : _GEN_1214; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1436 = 2'h1 == immu_state ? tlbl2_10_flag_v : _GEN_1215; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1437 = 2'h1 == immu_state ? tlbl2_11_flag_v : _GEN_1216; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1438 = 2'h1 == immu_state ? tlbl2_12_flag_v : _GEN_1217; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1439 = 2'h1 == immu_state ? tlbl2_13_flag_v : _GEN_1218; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1440 = 2'h1 == immu_state ? tlbl2_14_flag_v : _GEN_1219; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1441 = 2'h1 == immu_state ? tlbl2_15_flag_v : _GEN_1220; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1442 = 2'h1 == immu_state ? tlbl2_0_ppn : _GEN_1221; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1443 = 2'h1 == immu_state ? tlbl2_1_ppn : _GEN_1222; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1444 = 2'h1 == immu_state ? tlbl2_2_ppn : _GEN_1223; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1445 = 2'h1 == immu_state ? tlbl2_3_ppn : _GEN_1224; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1446 = 2'h1 == immu_state ? tlbl2_4_ppn : _GEN_1225; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1447 = 2'h1 == immu_state ? tlbl2_5_ppn : _GEN_1226; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1448 = 2'h1 == immu_state ? tlbl2_6_ppn : _GEN_1227; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1449 = 2'h1 == immu_state ? tlbl2_7_ppn : _GEN_1228; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1450 = 2'h1 == immu_state ? tlbl2_8_ppn : _GEN_1229; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1451 = 2'h1 == immu_state ? tlbl2_9_ppn : _GEN_1230; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1452 = 2'h1 == immu_state ? tlbl2_10_ppn : _GEN_1231; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1453 = 2'h1 == immu_state ? tlbl2_11_ppn : _GEN_1232; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1454 = 2'h1 == immu_state ? tlbl2_12_ppn : _GEN_1233; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1455 = 2'h1 == immu_state ? tlbl2_13_ppn : _GEN_1234; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1456 = 2'h1 == immu_state ? tlbl2_14_ppn : _GEN_1235; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1457 = 2'h1 == immu_state ? tlbl2_15_ppn : _GEN_1236; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1458 = 2'h1 == immu_state ? tlbl2_0_rmask : _GEN_1237; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1459 = 2'h1 == immu_state ? tlbl2_1_rmask : _GEN_1238; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1460 = 2'h1 == immu_state ? tlbl2_2_rmask : _GEN_1239; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1461 = 2'h1 == immu_state ? tlbl2_3_rmask : _GEN_1240; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1462 = 2'h1 == immu_state ? tlbl2_4_rmask : _GEN_1241; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1463 = 2'h1 == immu_state ? tlbl2_5_rmask : _GEN_1242; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1464 = 2'h1 == immu_state ? tlbl2_6_rmask : _GEN_1243; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1465 = 2'h1 == immu_state ? tlbl2_7_rmask : _GEN_1244; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1466 = 2'h1 == immu_state ? tlbl2_8_rmask : _GEN_1245; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1467 = 2'h1 == immu_state ? tlbl2_9_rmask : _GEN_1246; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1468 = 2'h1 == immu_state ? tlbl2_10_rmask : _GEN_1247; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1469 = 2'h1 == immu_state ? tlbl2_11_rmask : _GEN_1248; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1470 = 2'h1 == immu_state ? tlbl2_12_rmask : _GEN_1249; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1471 = 2'h1 == immu_state ? tlbl2_13_rmask : _GEN_1250; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1472 = 2'h1 == immu_state ? tlbl2_14_rmask : _GEN_1251; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1473 = 2'h1 == immu_state ? tlbl2_15_rmask : _GEN_1252; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [3:0] _GEN_1474 = 2'h1 == immu_state ? replace_index_value : _GEN_1265; // @[playground/src/cache/mmu/Tlb.scala 193:22 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _GEN_1488 = 2'h0 == immu_state ? itlb_flag_v : _GEN_1276; // @[playground/src/cache/mmu/Tlb.scala 193:22 75:22]
  wire [26:0] _GEN_1492 = 2'h0 == immu_state ? tlbl2_0_vpn : _GEN_1282; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1493 = 2'h0 == immu_state ? tlbl2_1_vpn : _GEN_1283; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1494 = 2'h0 == immu_state ? tlbl2_2_vpn : _GEN_1284; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1495 = 2'h0 == immu_state ? tlbl2_3_vpn : _GEN_1285; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1496 = 2'h0 == immu_state ? tlbl2_4_vpn : _GEN_1286; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1497 = 2'h0 == immu_state ? tlbl2_5_vpn : _GEN_1287; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1498 = 2'h0 == immu_state ? tlbl2_6_vpn : _GEN_1288; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1499 = 2'h0 == immu_state ? tlbl2_7_vpn : _GEN_1289; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1500 = 2'h0 == immu_state ? tlbl2_8_vpn : _GEN_1290; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1501 = 2'h0 == immu_state ? tlbl2_9_vpn : _GEN_1291; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1502 = 2'h0 == immu_state ? tlbl2_10_vpn : _GEN_1292; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1503 = 2'h0 == immu_state ? tlbl2_11_vpn : _GEN_1293; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1504 = 2'h0 == immu_state ? tlbl2_12_vpn : _GEN_1294; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1505 = 2'h0 == immu_state ? tlbl2_13_vpn : _GEN_1295; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1506 = 2'h0 == immu_state ? tlbl2_14_vpn : _GEN_1296; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [26:0] _GEN_1507 = 2'h0 == immu_state ? tlbl2_15_vpn : _GEN_1297; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1508 = 2'h0 == immu_state ? tlbl2_0_asid : _GEN_1298; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1509 = 2'h0 == immu_state ? tlbl2_1_asid : _GEN_1299; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1510 = 2'h0 == immu_state ? tlbl2_2_asid : _GEN_1300; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1511 = 2'h0 == immu_state ? tlbl2_3_asid : _GEN_1301; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1512 = 2'h0 == immu_state ? tlbl2_4_asid : _GEN_1302; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1513 = 2'h0 == immu_state ? tlbl2_5_asid : _GEN_1303; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1514 = 2'h0 == immu_state ? tlbl2_6_asid : _GEN_1304; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1515 = 2'h0 == immu_state ? tlbl2_7_asid : _GEN_1305; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1516 = 2'h0 == immu_state ? tlbl2_8_asid : _GEN_1306; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1517 = 2'h0 == immu_state ? tlbl2_9_asid : _GEN_1307; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1518 = 2'h0 == immu_state ? tlbl2_10_asid : _GEN_1308; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1519 = 2'h0 == immu_state ? tlbl2_11_asid : _GEN_1309; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1520 = 2'h0 == immu_state ? tlbl2_12_asid : _GEN_1310; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1521 = 2'h0 == immu_state ? tlbl2_13_asid : _GEN_1311; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1522 = 2'h0 == immu_state ? tlbl2_14_asid : _GEN_1312; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [15:0] _GEN_1523 = 2'h0 == immu_state ? tlbl2_15_asid : _GEN_1313; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1524 = 2'h0 == immu_state ? tlbl2_0_flag_d : _GEN_1314; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1525 = 2'h0 == immu_state ? tlbl2_1_flag_d : _GEN_1315; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1526 = 2'h0 == immu_state ? tlbl2_2_flag_d : _GEN_1316; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1527 = 2'h0 == immu_state ? tlbl2_3_flag_d : _GEN_1317; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1528 = 2'h0 == immu_state ? tlbl2_4_flag_d : _GEN_1318; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1529 = 2'h0 == immu_state ? tlbl2_5_flag_d : _GEN_1319; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1530 = 2'h0 == immu_state ? tlbl2_6_flag_d : _GEN_1320; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1531 = 2'h0 == immu_state ? tlbl2_7_flag_d : _GEN_1321; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1532 = 2'h0 == immu_state ? tlbl2_8_flag_d : _GEN_1322; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1533 = 2'h0 == immu_state ? tlbl2_9_flag_d : _GEN_1323; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1534 = 2'h0 == immu_state ? tlbl2_10_flag_d : _GEN_1324; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1535 = 2'h0 == immu_state ? tlbl2_11_flag_d : _GEN_1325; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1536 = 2'h0 == immu_state ? tlbl2_12_flag_d : _GEN_1326; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1537 = 2'h0 == immu_state ? tlbl2_13_flag_d : _GEN_1327; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1538 = 2'h0 == immu_state ? tlbl2_14_flag_d : _GEN_1328; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1539 = 2'h0 == immu_state ? tlbl2_15_flag_d : _GEN_1329; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1556 = 2'h0 == immu_state ? tlbl2_0_flag_g : _GEN_1346; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1557 = 2'h0 == immu_state ? tlbl2_1_flag_g : _GEN_1347; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1558 = 2'h0 == immu_state ? tlbl2_2_flag_g : _GEN_1348; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1559 = 2'h0 == immu_state ? tlbl2_3_flag_g : _GEN_1349; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1560 = 2'h0 == immu_state ? tlbl2_4_flag_g : _GEN_1350; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1561 = 2'h0 == immu_state ? tlbl2_5_flag_g : _GEN_1351; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1562 = 2'h0 == immu_state ? tlbl2_6_flag_g : _GEN_1352; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1563 = 2'h0 == immu_state ? tlbl2_7_flag_g : _GEN_1353; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1564 = 2'h0 == immu_state ? tlbl2_8_flag_g : _GEN_1354; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1565 = 2'h0 == immu_state ? tlbl2_9_flag_g : _GEN_1355; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1566 = 2'h0 == immu_state ? tlbl2_10_flag_g : _GEN_1356; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1567 = 2'h0 == immu_state ? tlbl2_11_flag_g : _GEN_1357; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1568 = 2'h0 == immu_state ? tlbl2_12_flag_g : _GEN_1358; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1569 = 2'h0 == immu_state ? tlbl2_13_flag_g : _GEN_1359; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1570 = 2'h0 == immu_state ? tlbl2_14_flag_g : _GEN_1360; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1571 = 2'h0 == immu_state ? tlbl2_15_flag_g : _GEN_1361; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1572 = 2'h0 == immu_state ? tlbl2_0_flag_u : _GEN_1362; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1573 = 2'h0 == immu_state ? tlbl2_1_flag_u : _GEN_1363; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1574 = 2'h0 == immu_state ? tlbl2_2_flag_u : _GEN_1364; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1575 = 2'h0 == immu_state ? tlbl2_3_flag_u : _GEN_1365; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1576 = 2'h0 == immu_state ? tlbl2_4_flag_u : _GEN_1366; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1577 = 2'h0 == immu_state ? tlbl2_5_flag_u : _GEN_1367; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1578 = 2'h0 == immu_state ? tlbl2_6_flag_u : _GEN_1368; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1579 = 2'h0 == immu_state ? tlbl2_7_flag_u : _GEN_1369; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1580 = 2'h0 == immu_state ? tlbl2_8_flag_u : _GEN_1370; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1581 = 2'h0 == immu_state ? tlbl2_9_flag_u : _GEN_1371; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1582 = 2'h0 == immu_state ? tlbl2_10_flag_u : _GEN_1372; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1583 = 2'h0 == immu_state ? tlbl2_11_flag_u : _GEN_1373; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1584 = 2'h0 == immu_state ? tlbl2_12_flag_u : _GEN_1374; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1585 = 2'h0 == immu_state ? tlbl2_13_flag_u : _GEN_1375; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1586 = 2'h0 == immu_state ? tlbl2_14_flag_u : _GEN_1376; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1587 = 2'h0 == immu_state ? tlbl2_15_flag_u : _GEN_1377; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1588 = 2'h0 == immu_state ? tlbl2_0_flag_x : _GEN_1378; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1589 = 2'h0 == immu_state ? tlbl2_1_flag_x : _GEN_1379; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1590 = 2'h0 == immu_state ? tlbl2_2_flag_x : _GEN_1380; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1591 = 2'h0 == immu_state ? tlbl2_3_flag_x : _GEN_1381; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1592 = 2'h0 == immu_state ? tlbl2_4_flag_x : _GEN_1382; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1593 = 2'h0 == immu_state ? tlbl2_5_flag_x : _GEN_1383; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1594 = 2'h0 == immu_state ? tlbl2_6_flag_x : _GEN_1384; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1595 = 2'h0 == immu_state ? tlbl2_7_flag_x : _GEN_1385; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1596 = 2'h0 == immu_state ? tlbl2_8_flag_x : _GEN_1386; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1597 = 2'h0 == immu_state ? tlbl2_9_flag_x : _GEN_1387; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1598 = 2'h0 == immu_state ? tlbl2_10_flag_x : _GEN_1388; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1599 = 2'h0 == immu_state ? tlbl2_11_flag_x : _GEN_1389; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1600 = 2'h0 == immu_state ? tlbl2_12_flag_x : _GEN_1390; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1601 = 2'h0 == immu_state ? tlbl2_13_flag_x : _GEN_1391; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1602 = 2'h0 == immu_state ? tlbl2_14_flag_x : _GEN_1392; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1603 = 2'h0 == immu_state ? tlbl2_15_flag_x : _GEN_1393; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1604 = 2'h0 == immu_state ? tlbl2_0_flag_w : _GEN_1394; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1605 = 2'h0 == immu_state ? tlbl2_1_flag_w : _GEN_1395; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1606 = 2'h0 == immu_state ? tlbl2_2_flag_w : _GEN_1396; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1607 = 2'h0 == immu_state ? tlbl2_3_flag_w : _GEN_1397; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1608 = 2'h0 == immu_state ? tlbl2_4_flag_w : _GEN_1398; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1609 = 2'h0 == immu_state ? tlbl2_5_flag_w : _GEN_1399; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1610 = 2'h0 == immu_state ? tlbl2_6_flag_w : _GEN_1400; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1611 = 2'h0 == immu_state ? tlbl2_7_flag_w : _GEN_1401; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1612 = 2'h0 == immu_state ? tlbl2_8_flag_w : _GEN_1402; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1613 = 2'h0 == immu_state ? tlbl2_9_flag_w : _GEN_1403; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1614 = 2'h0 == immu_state ? tlbl2_10_flag_w : _GEN_1404; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1615 = 2'h0 == immu_state ? tlbl2_11_flag_w : _GEN_1405; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1616 = 2'h0 == immu_state ? tlbl2_12_flag_w : _GEN_1406; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1617 = 2'h0 == immu_state ? tlbl2_13_flag_w : _GEN_1407; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1618 = 2'h0 == immu_state ? tlbl2_14_flag_w : _GEN_1408; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1619 = 2'h0 == immu_state ? tlbl2_15_flag_w : _GEN_1409; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1620 = 2'h0 == immu_state ? tlbl2_0_flag_r : _GEN_1410; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1621 = 2'h0 == immu_state ? tlbl2_1_flag_r : _GEN_1411; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1622 = 2'h0 == immu_state ? tlbl2_2_flag_r : _GEN_1412; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1623 = 2'h0 == immu_state ? tlbl2_3_flag_r : _GEN_1413; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1624 = 2'h0 == immu_state ? tlbl2_4_flag_r : _GEN_1414; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1625 = 2'h0 == immu_state ? tlbl2_5_flag_r : _GEN_1415; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1626 = 2'h0 == immu_state ? tlbl2_6_flag_r : _GEN_1416; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1627 = 2'h0 == immu_state ? tlbl2_7_flag_r : _GEN_1417; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1628 = 2'h0 == immu_state ? tlbl2_8_flag_r : _GEN_1418; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1629 = 2'h0 == immu_state ? tlbl2_9_flag_r : _GEN_1419; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1630 = 2'h0 == immu_state ? tlbl2_10_flag_r : _GEN_1420; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1631 = 2'h0 == immu_state ? tlbl2_11_flag_r : _GEN_1421; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1632 = 2'h0 == immu_state ? tlbl2_12_flag_r : _GEN_1422; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1633 = 2'h0 == immu_state ? tlbl2_13_flag_r : _GEN_1423; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1634 = 2'h0 == immu_state ? tlbl2_14_flag_r : _GEN_1424; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1635 = 2'h0 == immu_state ? tlbl2_15_flag_r : _GEN_1425; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1636 = 2'h0 == immu_state ? tlbl2_0_flag_v : _GEN_1426; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1637 = 2'h0 == immu_state ? tlbl2_1_flag_v : _GEN_1427; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1638 = 2'h0 == immu_state ? tlbl2_2_flag_v : _GEN_1428; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1639 = 2'h0 == immu_state ? tlbl2_3_flag_v : _GEN_1429; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1640 = 2'h0 == immu_state ? tlbl2_4_flag_v : _GEN_1430; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1641 = 2'h0 == immu_state ? tlbl2_5_flag_v : _GEN_1431; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1642 = 2'h0 == immu_state ? tlbl2_6_flag_v : _GEN_1432; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1643 = 2'h0 == immu_state ? tlbl2_7_flag_v : _GEN_1433; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1644 = 2'h0 == immu_state ? tlbl2_8_flag_v : _GEN_1434; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1645 = 2'h0 == immu_state ? tlbl2_9_flag_v : _GEN_1435; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1646 = 2'h0 == immu_state ? tlbl2_10_flag_v : _GEN_1436; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1647 = 2'h0 == immu_state ? tlbl2_11_flag_v : _GEN_1437; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1648 = 2'h0 == immu_state ? tlbl2_12_flag_v : _GEN_1438; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1649 = 2'h0 == immu_state ? tlbl2_13_flag_v : _GEN_1439; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1650 = 2'h0 == immu_state ? tlbl2_14_flag_v : _GEN_1440; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire  _GEN_1651 = 2'h0 == immu_state ? tlbl2_15_flag_v : _GEN_1441; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1652 = 2'h0 == immu_state ? tlbl2_0_ppn : _GEN_1442; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1653 = 2'h0 == immu_state ? tlbl2_1_ppn : _GEN_1443; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1654 = 2'h0 == immu_state ? tlbl2_2_ppn : _GEN_1444; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1655 = 2'h0 == immu_state ? tlbl2_3_ppn : _GEN_1445; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1656 = 2'h0 == immu_state ? tlbl2_4_ppn : _GEN_1446; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1657 = 2'h0 == immu_state ? tlbl2_5_ppn : _GEN_1447; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1658 = 2'h0 == immu_state ? tlbl2_6_ppn : _GEN_1448; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1659 = 2'h0 == immu_state ? tlbl2_7_ppn : _GEN_1449; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1660 = 2'h0 == immu_state ? tlbl2_8_ppn : _GEN_1450; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1661 = 2'h0 == immu_state ? tlbl2_9_ppn : _GEN_1451; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1662 = 2'h0 == immu_state ? tlbl2_10_ppn : _GEN_1452; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1663 = 2'h0 == immu_state ? tlbl2_11_ppn : _GEN_1453; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1664 = 2'h0 == immu_state ? tlbl2_12_ppn : _GEN_1454; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1665 = 2'h0 == immu_state ? tlbl2_13_ppn : _GEN_1455; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1666 = 2'h0 == immu_state ? tlbl2_14_ppn : _GEN_1456; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [19:0] _GEN_1667 = 2'h0 == immu_state ? tlbl2_15_ppn : _GEN_1457; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1668 = 2'h0 == immu_state ? tlbl2_0_rmask : _GEN_1458; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1669 = 2'h0 == immu_state ? tlbl2_1_rmask : _GEN_1459; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1670 = 2'h0 == immu_state ? tlbl2_2_rmask : _GEN_1460; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1671 = 2'h0 == immu_state ? tlbl2_3_rmask : _GEN_1461; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1672 = 2'h0 == immu_state ? tlbl2_4_rmask : _GEN_1462; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1673 = 2'h0 == immu_state ? tlbl2_5_rmask : _GEN_1463; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1674 = 2'h0 == immu_state ? tlbl2_6_rmask : _GEN_1464; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1675 = 2'h0 == immu_state ? tlbl2_7_rmask : _GEN_1465; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1676 = 2'h0 == immu_state ? tlbl2_8_rmask : _GEN_1466; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1677 = 2'h0 == immu_state ? tlbl2_9_rmask : _GEN_1467; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1678 = 2'h0 == immu_state ? tlbl2_10_rmask : _GEN_1468; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1679 = 2'h0 == immu_state ? tlbl2_11_rmask : _GEN_1469; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1680 = 2'h0 == immu_state ? tlbl2_12_rmask : _GEN_1470; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1681 = 2'h0 == immu_state ? tlbl2_13_rmask : _GEN_1471; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1682 = 2'h0 == immu_state ? tlbl2_14_rmask : _GEN_1472; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [17:0] _GEN_1683 = 2'h0 == immu_state ? tlbl2_15_rmask : _GEN_1473; // @[playground/src/cache/mmu/Tlb.scala 193:22 77:22]
  wire [3:0] _GEN_1684 = 2'h0 == immu_state ? replace_index_value : _GEN_1474; // @[playground/src/cache/mmu/Tlb.scala 193:22 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _T_17 = ~dtlb_flag_r; // @[playground/src/cache/mmu/Tlb.scala 285:22]
  wire  _T_22 = dtlb_flag_u & _T_4; // @[playground/src/cache/mmu/Tlb.scala 172:26]
  wire [1:0] _GEN_1686 = dtlb_flag_u & _T_4 ? 2'h3 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 172:42 174:23 107:76]
  wire  _GEN_1687 = dtlb_flag_u & _T_4 ? 1'h0 : 1'h1; // @[playground/src/cache/mmu/Tlb.scala 172:42 176:25 281:25]
  wire  _T_24 = ~dtlb_flag_u; // @[playground/src/cache/mmu/Tlb.scala 180:14]
  wire [1:0] _GEN_1689 = ~dtlb_flag_u ? 2'h3 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 180:28 182:23 107:76]
  wire  _GEN_1690 = ~dtlb_flag_u ? 1'h0 : 1'h1; // @[playground/src/cache/mmu/Tlb.scala 180:28 184:25 281:25]
  wire  _GEN_1691 = 2'h0 == io_csr_dmode & _T_24; // @[playground/src/cache/mmu/Tlb.scala 170:19 270:23]
  wire [1:0] _GEN_1692 = 2'h0 == io_csr_dmode ? _GEN_1689 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 170:19 107:76]
  wire  _GEN_1693 = 2'h0 == io_csr_dmode & _GEN_1690; // @[playground/src/cache/mmu/Tlb.scala 170:19 281:25]
  wire  _GEN_1694 = 2'h1 == io_csr_dmode ? _T_22 : _GEN_1691; // @[playground/src/cache/mmu/Tlb.scala 170:19]
  wire [1:0] _GEN_1695 = 2'h1 == io_csr_dmode ? _GEN_1686 : _GEN_1692; // @[playground/src/cache/mmu/Tlb.scala 170:19]
  wire  _GEN_1696 = 2'h1 == io_csr_dmode ? _GEN_1687 : _GEN_1693; // @[playground/src/cache/mmu/Tlb.scala 170:19]
  wire  _GEN_1697 = ~dtlb_flag_r & ~dtlb_flag_x | _GEN_1694; // @[playground/src/cache/mmu/Tlb.scala 285:52 286:31]
  wire [1:0] _GEN_1698 = ~dtlb_flag_r & ~dtlb_flag_x ? 2'h3 : _GEN_1695; // @[playground/src/cache/mmu/Tlb.scala 285:52 287:31]
  wire  _GEN_1699 = ~dtlb_flag_r & ~dtlb_flag_x ? 1'h0 : _GEN_1696; // @[playground/src/cache/mmu/Tlb.scala 281:25 285:52]
  wire  _GEN_1712 = _T_17 | _GEN_1694; // @[playground/src/cache/mmu/Tlb.scala 292:36 293:31]
  wire [1:0] _GEN_1713 = _T_17 ? 2'h3 : _GEN_1695; // @[playground/src/cache/mmu/Tlb.scala 292:36 294:31]
  wire  _GEN_1714 = _T_17 ? 1'h0 : _GEN_1696; // @[playground/src/cache/mmu/Tlb.scala 281:25 292:36]
  wire  _GEN_1715 = mstatus_mxr ? _GEN_1697 : _GEN_1712; // @[playground/src/cache/mmu/Tlb.scala 284:25]
  wire [1:0] _GEN_1716 = mstatus_mxr ? _GEN_1698 : _GEN_1713; // @[playground/src/cache/mmu/Tlb.scala 284:25]
  wire  _GEN_1717 = mstatus_mxr ? _GEN_1699 : _GEN_1714; // @[playground/src/cache/mmu/Tlb.scala 284:25]
  wire  _GEN_1730 = ~dtlb_flag_w | _GEN_1694; // @[playground/src/cache/mmu/Tlb.scala 305:36 306:31]
  wire [1:0] _GEN_1731 = ~dtlb_flag_w ? 2'h3 : _GEN_1695; // @[playground/src/cache/mmu/Tlb.scala 305:36 307:31]
  wire  _GEN_1732 = ~dtlb_flag_w ? 1'h0 : _GEN_1696; // @[playground/src/cache/mmu/Tlb.scala 281:25 305:36]
  wire  _GEN_1733 = ~dtlb_flag_d | _GEN_1730; // @[playground/src/cache/mmu/Tlb.scala 301:34 302:29]
  wire [1:0] _GEN_1734 = ~dtlb_flag_d ? 2'h3 : _GEN_1731; // @[playground/src/cache/mmu/Tlb.scala 301:34 303:29]
  wire  _GEN_1735 = ~dtlb_flag_d ? 1'h0 : _GEN_1732; // @[playground/src/cache/mmu/Tlb.scala 281:25 301:34]
  wire  _GEN_1736 = 2'h2 == io_dcache_access_type & _GEN_1733; // @[playground/src/cache/mmu/Tlb.scala 270:23 282:41]
  wire [1:0] _GEN_1737 = 2'h2 == io_dcache_access_type ? _GEN_1734 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 282:41 107:76]
  wire  _GEN_1738 = 2'h2 == io_dcache_access_type & _GEN_1735; // @[playground/src/cache/mmu/Tlb.scala 281:25 282:41]
  wire  _GEN_1739 = 2'h1 == io_dcache_access_type ? _GEN_1715 : _GEN_1736; // @[playground/src/cache/mmu/Tlb.scala 282:41]
  wire [1:0] _GEN_1740 = 2'h1 == io_dcache_access_type ? _GEN_1716 : _GEN_1737; // @[playground/src/cache/mmu/Tlb.scala 282:41]
  wire  _GEN_1741 = 2'h1 == io_dcache_access_type ? _GEN_1717 : _GEN_1738; // @[playground/src/cache/mmu/Tlb.scala 282:41]
  wire  _GEN_1742 = dtlbl1_hit & _GEN_1741; // @[playground/src/cache/mmu/Tlb.scala 135:26 274:32]
  wire  _GEN_1743 = dtlbl1_hit & _GEN_1739; // @[playground/src/cache/mmu/Tlb.scala 270:23 274:32]
  wire [1:0] _GEN_1744 = dtlbl1_hit ? _GEN_1740 : 2'h1; // @[playground/src/cache/mmu/Tlb.scala 274:32 315:22]
  wire  _GEN_1745 = ~dvm_enabled | _GEN_1742; // @[playground/src/cache/mmu/Tlb.scala 272:28 273:25]
  wire  _GEN_1750 = io_dcache_en & _GEN_1745; // @[playground/src/cache/mmu/Tlb.scala 135:26 268:26]
  wire [3:0] _dtlb_T = dl2_hit_vec_14 ? 4'he : 4'hf; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_1 = dl2_hit_vec_13 ? 4'hd : _dtlb_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_2 = dl2_hit_vec_12 ? 4'hc : _dtlb_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_3 = dl2_hit_vec_11 ? 4'hb : _dtlb_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_4 = dl2_hit_vec_10 ? 4'ha : _dtlb_T_3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_5 = dl2_hit_vec_9 ? 4'h9 : _dtlb_T_4; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_6 = dl2_hit_vec_8 ? 4'h8 : _dtlb_T_5; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_7 = dl2_hit_vec_7 ? 4'h7 : _dtlb_T_6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_8 = dl2_hit_vec_6 ? 4'h6 : _dtlb_T_7; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_9 = dl2_hit_vec_5 ? 4'h5 : _dtlb_T_8; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_10 = dl2_hit_vec_4 ? 4'h4 : _dtlb_T_9; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_11 = dl2_hit_vec_3 ? 4'h3 : _dtlb_T_10; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_12 = dl2_hit_vec_2 ? 4'h2 : _dtlb_T_11; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_13 = dl2_hit_vec_1 ? 4'h1 : _dtlb_T_12; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _dtlb_T_14 = dl2_hit_vec_0 ? 4'h0 : _dtlb_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [26:0] _GEN_1753 = 4'h1 == _dtlb_T_14 ? tlbl2_1_vpn : tlbl2_0_vpn; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1754 = 4'h2 == _dtlb_T_14 ? tlbl2_2_vpn : _GEN_1753; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1755 = 4'h3 == _dtlb_T_14 ? tlbl2_3_vpn : _GEN_1754; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1756 = 4'h4 == _dtlb_T_14 ? tlbl2_4_vpn : _GEN_1755; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1757 = 4'h5 == _dtlb_T_14 ? tlbl2_5_vpn : _GEN_1756; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1758 = 4'h6 == _dtlb_T_14 ? tlbl2_6_vpn : _GEN_1757; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1759 = 4'h7 == _dtlb_T_14 ? tlbl2_7_vpn : _GEN_1758; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1760 = 4'h8 == _dtlb_T_14 ? tlbl2_8_vpn : _GEN_1759; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1761 = 4'h9 == _dtlb_T_14 ? tlbl2_9_vpn : _GEN_1760; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1762 = 4'ha == _dtlb_T_14 ? tlbl2_10_vpn : _GEN_1761; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1763 = 4'hb == _dtlb_T_14 ? tlbl2_11_vpn : _GEN_1762; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1764 = 4'hc == _dtlb_T_14 ? tlbl2_12_vpn : _GEN_1763; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1765 = 4'hd == _dtlb_T_14 ? tlbl2_13_vpn : _GEN_1764; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1766 = 4'he == _dtlb_T_14 ? tlbl2_14_vpn : _GEN_1765; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [26:0] _GEN_1767 = 4'hf == _dtlb_T_14 ? tlbl2_15_vpn : _GEN_1766; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1769 = 4'h1 == _dtlb_T_14 ? tlbl2_1_asid : tlbl2_0_asid; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1770 = 4'h2 == _dtlb_T_14 ? tlbl2_2_asid : _GEN_1769; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1771 = 4'h3 == _dtlb_T_14 ? tlbl2_3_asid : _GEN_1770; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1772 = 4'h4 == _dtlb_T_14 ? tlbl2_4_asid : _GEN_1771; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1773 = 4'h5 == _dtlb_T_14 ? tlbl2_5_asid : _GEN_1772; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1774 = 4'h6 == _dtlb_T_14 ? tlbl2_6_asid : _GEN_1773; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1775 = 4'h7 == _dtlb_T_14 ? tlbl2_7_asid : _GEN_1774; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1776 = 4'h8 == _dtlb_T_14 ? tlbl2_8_asid : _GEN_1775; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1777 = 4'h9 == _dtlb_T_14 ? tlbl2_9_asid : _GEN_1776; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1778 = 4'ha == _dtlb_T_14 ? tlbl2_10_asid : _GEN_1777; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1779 = 4'hb == _dtlb_T_14 ? tlbl2_11_asid : _GEN_1778; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1780 = 4'hc == _dtlb_T_14 ? tlbl2_12_asid : _GEN_1779; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1781 = 4'hd == _dtlb_T_14 ? tlbl2_13_asid : _GEN_1780; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1782 = 4'he == _dtlb_T_14 ? tlbl2_14_asid : _GEN_1781; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [15:0] _GEN_1783 = 4'hf == _dtlb_T_14 ? tlbl2_15_asid : _GEN_1782; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1785 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_d : tlbl2_0_flag_d; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1786 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_d : _GEN_1785; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1787 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_d : _GEN_1786; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1788 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_d : _GEN_1787; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1789 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_d : _GEN_1788; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1790 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_d : _GEN_1789; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1791 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_d : _GEN_1790; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1792 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_d : _GEN_1791; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1793 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_d : _GEN_1792; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1794 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_d : _GEN_1793; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1795 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_d : _GEN_1794; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1796 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_d : _GEN_1795; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1797 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_d : _GEN_1796; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1798 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_d : _GEN_1797; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1799 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_d : _GEN_1798; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1817 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_g : tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1818 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_g : _GEN_1817; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1819 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_g : _GEN_1818; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1820 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_g : _GEN_1819; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1821 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_g : _GEN_1820; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1822 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_g : _GEN_1821; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1823 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_g : _GEN_1822; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1824 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_g : _GEN_1823; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1825 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_g : _GEN_1824; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1826 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_g : _GEN_1825; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1827 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_g : _GEN_1826; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1828 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_g : _GEN_1827; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1829 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_g : _GEN_1828; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1830 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_g : _GEN_1829; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1831 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_g : _GEN_1830; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1833 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_u : tlbl2_0_flag_u; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1834 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_u : _GEN_1833; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1835 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_u : _GEN_1834; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1836 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_u : _GEN_1835; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1837 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_u : _GEN_1836; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1838 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_u : _GEN_1837; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1839 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_u : _GEN_1838; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1840 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_u : _GEN_1839; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1841 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_u : _GEN_1840; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1842 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_u : _GEN_1841; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1843 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_u : _GEN_1842; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1844 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_u : _GEN_1843; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1845 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_u : _GEN_1844; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1846 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_u : _GEN_1845; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1847 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_u : _GEN_1846; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1849 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_x : tlbl2_0_flag_x; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1850 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_x : _GEN_1849; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1851 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_x : _GEN_1850; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1852 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_x : _GEN_1851; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1853 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_x : _GEN_1852; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1854 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_x : _GEN_1853; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1855 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_x : _GEN_1854; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1856 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_x : _GEN_1855; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1857 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_x : _GEN_1856; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1858 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_x : _GEN_1857; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1859 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_x : _GEN_1858; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1860 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_x : _GEN_1859; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1861 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_x : _GEN_1860; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1862 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_x : _GEN_1861; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1863 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_x : _GEN_1862; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1865 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_w : tlbl2_0_flag_w; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1866 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_w : _GEN_1865; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1867 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_w : _GEN_1866; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1868 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_w : _GEN_1867; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1869 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_w : _GEN_1868; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1870 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_w : _GEN_1869; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1871 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_w : _GEN_1870; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1872 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_w : _GEN_1871; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1873 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_w : _GEN_1872; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1874 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_w : _GEN_1873; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1875 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_w : _GEN_1874; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1876 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_w : _GEN_1875; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1877 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_w : _GEN_1876; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1878 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_w : _GEN_1877; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1879 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_w : _GEN_1878; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1881 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_r : tlbl2_0_flag_r; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1882 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_r : _GEN_1881; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1883 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_r : _GEN_1882; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1884 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_r : _GEN_1883; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1885 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_r : _GEN_1884; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1886 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_r : _GEN_1885; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1887 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_r : _GEN_1886; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1888 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_r : _GEN_1887; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1889 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_r : _GEN_1888; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1890 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_r : _GEN_1889; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1891 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_r : _GEN_1890; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1892 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_r : _GEN_1891; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1893 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_r : _GEN_1892; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1894 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_r : _GEN_1893; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1895 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_r : _GEN_1894; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1897 = 4'h1 == _dtlb_T_14 ? tlbl2_1_flag_v : tlbl2_0_flag_v; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1898 = 4'h2 == _dtlb_T_14 ? tlbl2_2_flag_v : _GEN_1897; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1899 = 4'h3 == _dtlb_T_14 ? tlbl2_3_flag_v : _GEN_1898; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1900 = 4'h4 == _dtlb_T_14 ? tlbl2_4_flag_v : _GEN_1899; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1901 = 4'h5 == _dtlb_T_14 ? tlbl2_5_flag_v : _GEN_1900; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1902 = 4'h6 == _dtlb_T_14 ? tlbl2_6_flag_v : _GEN_1901; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1903 = 4'h7 == _dtlb_T_14 ? tlbl2_7_flag_v : _GEN_1902; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1904 = 4'h8 == _dtlb_T_14 ? tlbl2_8_flag_v : _GEN_1903; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1905 = 4'h9 == _dtlb_T_14 ? tlbl2_9_flag_v : _GEN_1904; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1906 = 4'ha == _dtlb_T_14 ? tlbl2_10_flag_v : _GEN_1905; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1907 = 4'hb == _dtlb_T_14 ? tlbl2_11_flag_v : _GEN_1906; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1908 = 4'hc == _dtlb_T_14 ? tlbl2_12_flag_v : _GEN_1907; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1909 = 4'hd == _dtlb_T_14 ? tlbl2_13_flag_v : _GEN_1908; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1910 = 4'he == _dtlb_T_14 ? tlbl2_14_flag_v : _GEN_1909; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire  _GEN_1911 = 4'hf == _dtlb_T_14 ? tlbl2_15_flag_v : _GEN_1910; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1913 = 4'h1 == _dtlb_T_14 ? tlbl2_1_ppn : tlbl2_0_ppn; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1914 = 4'h2 == _dtlb_T_14 ? tlbl2_2_ppn : _GEN_1913; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1915 = 4'h3 == _dtlb_T_14 ? tlbl2_3_ppn : _GEN_1914; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1916 = 4'h4 == _dtlb_T_14 ? tlbl2_4_ppn : _GEN_1915; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1917 = 4'h5 == _dtlb_T_14 ? tlbl2_5_ppn : _GEN_1916; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1918 = 4'h6 == _dtlb_T_14 ? tlbl2_6_ppn : _GEN_1917; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1919 = 4'h7 == _dtlb_T_14 ? tlbl2_7_ppn : _GEN_1918; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1920 = 4'h8 == _dtlb_T_14 ? tlbl2_8_ppn : _GEN_1919; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1921 = 4'h9 == _dtlb_T_14 ? tlbl2_9_ppn : _GEN_1920; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1922 = 4'ha == _dtlb_T_14 ? tlbl2_10_ppn : _GEN_1921; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1923 = 4'hb == _dtlb_T_14 ? tlbl2_11_ppn : _GEN_1922; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1924 = 4'hc == _dtlb_T_14 ? tlbl2_12_ppn : _GEN_1923; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1925 = 4'hd == _dtlb_T_14 ? tlbl2_13_ppn : _GEN_1924; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1926 = 4'he == _dtlb_T_14 ? tlbl2_14_ppn : _GEN_1925; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [19:0] _GEN_1927 = 4'hf == _dtlb_T_14 ? tlbl2_15_ppn : _GEN_1926; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1929 = 4'h1 == _dtlb_T_14 ? tlbl2_1_rmask : tlbl2_0_rmask; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1930 = 4'h2 == _dtlb_T_14 ? tlbl2_2_rmask : _GEN_1929; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1931 = 4'h3 == _dtlb_T_14 ? tlbl2_3_rmask : _GEN_1930; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1932 = 4'h4 == _dtlb_T_14 ? tlbl2_4_rmask : _GEN_1931; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1933 = 4'h5 == _dtlb_T_14 ? tlbl2_5_rmask : _GEN_1932; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1934 = 4'h6 == _dtlb_T_14 ? tlbl2_6_rmask : _GEN_1933; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1935 = 4'h7 == _dtlb_T_14 ? tlbl2_7_rmask : _GEN_1934; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1936 = 4'h8 == _dtlb_T_14 ? tlbl2_8_rmask : _GEN_1935; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1937 = 4'h9 == _dtlb_T_14 ? tlbl2_9_rmask : _GEN_1936; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1938 = 4'ha == _dtlb_T_14 ? tlbl2_10_rmask : _GEN_1937; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1939 = 4'hb == _dtlb_T_14 ? tlbl2_11_rmask : _GEN_1938; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1940 = 4'hc == _dtlb_T_14 ? tlbl2_12_rmask : _GEN_1939; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1941 = 4'hd == _dtlb_T_14 ? tlbl2_13_rmask : _GEN_1940; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1942 = 4'he == _dtlb_T_14 ? tlbl2_14_rmask : _GEN_1941; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [17:0] _GEN_1943 = 4'hf == _dtlb_T_14 ? tlbl2_15_rmask : _GEN_1942; // @[playground/src/cache/mmu/Tlb.scala 322:{20,20}]
  wire [1:0] _GEN_1944 = ~choose_icache & io_dcache_ptw_vpn_ready ? 2'h2 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 325:57 326:22 107:76]
  wire  _GEN_1955 = |_T_40 ? _GEN_1911 : dtlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 320:36 322:20 76:22]
  wire [26:0] _GEN_1959 = 4'h0 == replace_index_value ? dvpn : _GEN_1492; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1960 = 4'h1 == replace_index_value ? dvpn : _GEN_1493; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1961 = 4'h2 == replace_index_value ? dvpn : _GEN_1494; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1962 = 4'h3 == replace_index_value ? dvpn : _GEN_1495; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1963 = 4'h4 == replace_index_value ? dvpn : _GEN_1496; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1964 = 4'h5 == replace_index_value ? dvpn : _GEN_1497; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1965 = 4'h6 == replace_index_value ? dvpn : _GEN_1498; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1966 = 4'h7 == replace_index_value ? dvpn : _GEN_1499; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1967 = 4'h8 == replace_index_value ? dvpn : _GEN_1500; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1968 = 4'h9 == replace_index_value ? dvpn : _GEN_1501; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1969 = 4'ha == replace_index_value ? dvpn : _GEN_1502; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1970 = 4'hb == replace_index_value ? dvpn : _GEN_1503; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1971 = 4'hc == replace_index_value ? dvpn : _GEN_1504; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1972 = 4'hd == replace_index_value ? dvpn : _GEN_1505; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1973 = 4'he == replace_index_value ? dvpn : _GEN_1506; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [26:0] _GEN_1974 = 4'hf == replace_index_value ? dvpn : _GEN_1507; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1975 = 4'h0 == replace_index_value ? satp_asid : _GEN_1508; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1976 = 4'h1 == replace_index_value ? satp_asid : _GEN_1509; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1977 = 4'h2 == replace_index_value ? satp_asid : _GEN_1510; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1978 = 4'h3 == replace_index_value ? satp_asid : _GEN_1511; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1979 = 4'h4 == replace_index_value ? satp_asid : _GEN_1512; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1980 = 4'h5 == replace_index_value ? satp_asid : _GEN_1513; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1981 = 4'h6 == replace_index_value ? satp_asid : _GEN_1514; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1982 = 4'h7 == replace_index_value ? satp_asid : _GEN_1515; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1983 = 4'h8 == replace_index_value ? satp_asid : _GEN_1516; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1984 = 4'h9 == replace_index_value ? satp_asid : _GEN_1517; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1985 = 4'ha == replace_index_value ? satp_asid : _GEN_1518; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1986 = 4'hb == replace_index_value ? satp_asid : _GEN_1519; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1987 = 4'hc == replace_index_value ? satp_asid : _GEN_1520; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1988 = 4'hd == replace_index_value ? satp_asid : _GEN_1521; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1989 = 4'he == replace_index_value ? satp_asid : _GEN_1522; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [15:0] _GEN_1990 = 4'hf == replace_index_value ? satp_asid : _GEN_1523; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1991 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1524; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1992 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1525; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1993 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1526; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1994 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1527; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1995 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1528; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1996 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1529; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1997 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1530; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1998 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1531; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_1999 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1532; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2000 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1533; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2001 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1534; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2002 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1535; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2003 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1536; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2004 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1537; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2005 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1538; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2006 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_d : _GEN_1539; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2023 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1556; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2024 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1557; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2025 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1558; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2026 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1559; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2027 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1560; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2028 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1561; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2029 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1562; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2030 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1563; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2031 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1564; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2032 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1565; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2033 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1566; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2034 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1567; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2035 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1568; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2036 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1569; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2037 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1570; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2038 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_g : _GEN_1571; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2039 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1572; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2040 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1573; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2041 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1574; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2042 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1575; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2043 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1576; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2044 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1577; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2045 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1578; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2046 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1579; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2047 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1580; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2048 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1581; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2049 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1582; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2050 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1583; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2051 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1584; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2052 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1585; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2053 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1586; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2054 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_u : _GEN_1587; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2055 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1588; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2056 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1589; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2057 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1590; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2058 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1591; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2059 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1592; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2060 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1593; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2061 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1594; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2062 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1595; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2063 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1596; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2064 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1597; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2065 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1598; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2066 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1599; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2067 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1600; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2068 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1601; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2069 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1602; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2070 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_x : _GEN_1603; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2071 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1604; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2072 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1605; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2073 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1606; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2074 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1607; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2075 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1608; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2076 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1609; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2077 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1610; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2078 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1611; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2079 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1612; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2080 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1613; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2081 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1614; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2082 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1615; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2083 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1616; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2084 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1617; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2085 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1618; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2086 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_w : _GEN_1619; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2087 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1620; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2088 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1621; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2089 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1622; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2090 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1623; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2091 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1624; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2092 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1625; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2093 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1626; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2094 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1627; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2095 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1628; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2096 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1629; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2097 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1630; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2098 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1631; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2099 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1632; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2100 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1633; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2101 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1634; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2102 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_r : _GEN_1635; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2103 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1636; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2104 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1637; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2105 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1638; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2106 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1639; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2107 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1640; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2108 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1641; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2109 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1642; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2110 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1643; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2111 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1644; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2112 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1645; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2113 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1646; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2114 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1647; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2115 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1648; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2116 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1649; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2117 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1650; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2118 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_flag_v : _GEN_1651; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2119 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1652; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2120 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1653; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2121 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1654; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2122 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1655; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2123 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1656; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2124 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1657; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2125 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1658; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2126 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1659; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2127 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1660; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2128 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1661; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2129 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1662; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2130 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1663; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2131 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1664; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2132 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1665; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2133 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1666; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [19:0] _GEN_2134 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_entry_ppn : _GEN_1667; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2135 = 4'h0 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1668; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2136 = 4'h1 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1669; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2137 = 4'h2 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1670; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2138 = 4'h3 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1671; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2139 = 4'h4 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1672; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2140 = 4'h5 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1673; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2141 = 4'h6 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1674; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2142 = 4'h7 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1675; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2143 = 4'h8 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1676; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2144 = 4'h9 == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1677; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2145 = 4'ha == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1678; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2146 = 4'hb == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1679; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2147 = 4'hc == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1680; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2148 = 4'hd == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1681; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2149 = 4'he == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1682; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire [17:0] _GEN_2150 = 4'hf == replace_index_value ? io_dcache_ptw_pte_bits_rmask : _GEN_1683; // @[playground/src/cache/mmu/Tlb.scala 347:{38,38}]
  wire  _GEN_2151 = io_dcache_ptw_pte_bits_page_fault | dpage_fault; // @[playground/src/cache/mmu/Tlb.scala 336:55 337:23 113:30]
  wire [26:0] _GEN_2152 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1492 : _GEN_1959; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2153 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1493 : _GEN_1960; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2154 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1494 : _GEN_1961; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2155 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1495 : _GEN_1962; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2156 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1496 : _GEN_1963; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2157 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1497 : _GEN_1964; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2158 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1498 : _GEN_1965; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2159 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1499 : _GEN_1966; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2160 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1500 : _GEN_1967; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2161 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1501 : _GEN_1968; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2162 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1502 : _GEN_1969; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2163 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1503 : _GEN_1970; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2164 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1504 : _GEN_1971; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2165 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1505 : _GEN_1972; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2166 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1506 : _GEN_1973; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2167 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1507 : _GEN_1974; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2168 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1508 : _GEN_1975; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2169 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1509 : _GEN_1976; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2170 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1510 : _GEN_1977; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2171 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1511 : _GEN_1978; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2172 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1512 : _GEN_1979; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2173 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1513 : _GEN_1980; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2174 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1514 : _GEN_1981; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2175 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1515 : _GEN_1982; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2176 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1516 : _GEN_1983; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2177 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1517 : _GEN_1984; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2178 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1518 : _GEN_1985; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2179 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1519 : _GEN_1986; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2180 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1520 : _GEN_1987; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2181 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1521 : _GEN_1988; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2182 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1522 : _GEN_1989; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [15:0] _GEN_2183 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1523 : _GEN_1990; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2184 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1524 : _GEN_1991; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2185 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1525 : _GEN_1992; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2186 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1526 : _GEN_1993; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2187 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1527 : _GEN_1994; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2188 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1528 : _GEN_1995; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2189 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1529 : _GEN_1996; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2190 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1530 : _GEN_1997; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2191 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1531 : _GEN_1998; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2192 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1532 : _GEN_1999; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2193 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1533 : _GEN_2000; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2194 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1534 : _GEN_2001; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2195 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1535 : _GEN_2002; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2196 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1536 : _GEN_2003; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2197 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1537 : _GEN_2004; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2198 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1538 : _GEN_2005; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2199 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1539 : _GEN_2006; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2216 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1556 : _GEN_2023; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2217 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1557 : _GEN_2024; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2218 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1558 : _GEN_2025; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2219 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1559 : _GEN_2026; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2220 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1560 : _GEN_2027; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2221 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1561 : _GEN_2028; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2222 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1562 : _GEN_2029; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2223 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1563 : _GEN_2030; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2224 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1564 : _GEN_2031; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2225 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1565 : _GEN_2032; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2226 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1566 : _GEN_2033; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2227 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1567 : _GEN_2034; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2228 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1568 : _GEN_2035; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2229 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1569 : _GEN_2036; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2230 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1570 : _GEN_2037; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2231 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1571 : _GEN_2038; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2232 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1572 : _GEN_2039; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2233 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1573 : _GEN_2040; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2234 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1574 : _GEN_2041; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2235 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1575 : _GEN_2042; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2236 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1576 : _GEN_2043; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2237 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1577 : _GEN_2044; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2238 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1578 : _GEN_2045; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2239 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1579 : _GEN_2046; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2240 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1580 : _GEN_2047; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2241 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1581 : _GEN_2048; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2242 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1582 : _GEN_2049; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2243 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1583 : _GEN_2050; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2244 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1584 : _GEN_2051; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2245 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1585 : _GEN_2052; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2246 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1586 : _GEN_2053; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2247 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1587 : _GEN_2054; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2248 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1588 : _GEN_2055; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2249 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1589 : _GEN_2056; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2250 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1590 : _GEN_2057; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2251 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1591 : _GEN_2058; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2252 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1592 : _GEN_2059; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2253 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1593 : _GEN_2060; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2254 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1594 : _GEN_2061; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2255 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1595 : _GEN_2062; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2256 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1596 : _GEN_2063; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2257 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1597 : _GEN_2064; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2258 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1598 : _GEN_2065; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2259 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1599 : _GEN_2066; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2260 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1600 : _GEN_2067; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2261 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1601 : _GEN_2068; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2262 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1602 : _GEN_2069; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2263 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1603 : _GEN_2070; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2264 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1604 : _GEN_2071; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2265 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1605 : _GEN_2072; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2266 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1606 : _GEN_2073; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2267 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1607 : _GEN_2074; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2268 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1608 : _GEN_2075; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2269 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1609 : _GEN_2076; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2270 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1610 : _GEN_2077; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2271 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1611 : _GEN_2078; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2272 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1612 : _GEN_2079; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2273 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1613 : _GEN_2080; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2274 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1614 : _GEN_2081; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2275 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1615 : _GEN_2082; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2276 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1616 : _GEN_2083; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2277 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1617 : _GEN_2084; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2278 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1618 : _GEN_2085; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2279 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1619 : _GEN_2086; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2280 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1620 : _GEN_2087; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2281 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1621 : _GEN_2088; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2282 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1622 : _GEN_2089; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2283 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1623 : _GEN_2090; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2284 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1624 : _GEN_2091; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2285 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1625 : _GEN_2092; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2286 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1626 : _GEN_2093; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2287 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1627 : _GEN_2094; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2288 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1628 : _GEN_2095; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2289 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1629 : _GEN_2096; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2290 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1630 : _GEN_2097; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2291 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1631 : _GEN_2098; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2292 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1632 : _GEN_2099; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2293 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1633 : _GEN_2100; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2294 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1634 : _GEN_2101; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2295 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1635 : _GEN_2102; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2296 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1636 : _GEN_2103; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2297 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1637 : _GEN_2104; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2298 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1638 : _GEN_2105; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2299 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1639 : _GEN_2106; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2300 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1640 : _GEN_2107; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2301 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1641 : _GEN_2108; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2302 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1642 : _GEN_2109; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2303 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1643 : _GEN_2110; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2304 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1644 : _GEN_2111; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2305 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1645 : _GEN_2112; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2306 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1646 : _GEN_2113; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2307 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1647 : _GEN_2114; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2308 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1648 : _GEN_2115; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2309 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1649 : _GEN_2116; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2310 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1650 : _GEN_2117; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire  _GEN_2311 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1651 : _GEN_2118; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2312 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1652 : _GEN_2119; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2313 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1653 : _GEN_2120; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2314 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1654 : _GEN_2121; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2315 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1655 : _GEN_2122; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2316 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1656 : _GEN_2123; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2317 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1657 : _GEN_2124; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2318 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1658 : _GEN_2125; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2319 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1659 : _GEN_2126; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2320 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1660 : _GEN_2127; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2321 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1661 : _GEN_2128; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2322 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1662 : _GEN_2129; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2323 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1663 : _GEN_2130; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2324 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1664 : _GEN_2131; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2325 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1665 : _GEN_2132; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2326 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1666 : _GEN_2133; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [19:0] _GEN_2327 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1667 : _GEN_2134; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2328 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1668 : _GEN_2135; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2329 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1669 : _GEN_2136; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2330 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1670 : _GEN_2137; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2331 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1671 : _GEN_2138; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2332 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1672 : _GEN_2139; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2333 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1673 : _GEN_2140; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2334 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1674 : _GEN_2141; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2335 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1675 : _GEN_2142; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2336 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1676 : _GEN_2143; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2337 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1677 : _GEN_2144; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2338 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1678 : _GEN_2145; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2339 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1679 : _GEN_2146; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2340 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1680 : _GEN_2147; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2341 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1681 : _GEN_2148; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2342 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1682 : _GEN_2149; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [17:0] _GEN_2343 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1683 : _GEN_2150; // @[playground/src/cache/mmu/Tlb.scala 336:55]
  wire [26:0] _GEN_2344 = io_dcache_ptw_pte_bits_page_fault ? dtlb_vpn : dvpn; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire [15:0] _GEN_2345 = io_dcache_ptw_pte_bits_page_fault ? dtlb_asid : satp_asid; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2346 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_d : io_dcache_ptw_pte_bits_entry_flag_d; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2348 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_g : io_dcache_ptw_pte_bits_entry_flag_g; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2349 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_u : io_dcache_ptw_pte_bits_entry_flag_u; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2350 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_x : io_dcache_ptw_pte_bits_entry_flag_x; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2351 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_w : io_dcache_ptw_pte_bits_entry_flag_w; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2352 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_r : io_dcache_ptw_pte_bits_entry_flag_r; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire  _GEN_2353 = io_dcache_ptw_pte_bits_page_fault ? dtlb_flag_v : io_dcache_ptw_pte_bits_entry_flag_v; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire [19:0] _GEN_2354 = io_dcache_ptw_pte_bits_page_fault ? dtlb_ppn : io_dcache_ptw_pte_bits_entry_ppn; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire [17:0] _GEN_2355 = io_dcache_ptw_pte_bits_page_fault ? dtlb_rmask : io_dcache_ptw_pte_bits_rmask; // @[playground/src/cache/mmu/Tlb.scala 336:55 76:22 348:38]
  wire [3:0] _GEN_2356 = io_dcache_ptw_pte_bits_page_fault ? _GEN_1684 : _value_T_1; // @[playground/src/cache/mmu/Tlb.scala 336:55 src/main/scala/chisel3/util/Counter.scala 77:15]
  wire [1:0] _GEN_2565 = io_dcache_ptw_pte_valid ? _GEN_429 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 332:37 107:76]
  wire  _GEN_2566 = io_dcache_ptw_pte_valid ? _GEN_2151 : dpage_fault; // @[playground/src/cache/mmu/Tlb.scala 113:30 332:37]
  wire [26:0] _GEN_2567 = io_dcache_ptw_pte_valid ? _GEN_2152 : _GEN_1492; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2568 = io_dcache_ptw_pte_valid ? _GEN_2153 : _GEN_1493; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2569 = io_dcache_ptw_pte_valid ? _GEN_2154 : _GEN_1494; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2570 = io_dcache_ptw_pte_valid ? _GEN_2155 : _GEN_1495; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2571 = io_dcache_ptw_pte_valid ? _GEN_2156 : _GEN_1496; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2572 = io_dcache_ptw_pte_valid ? _GEN_2157 : _GEN_1497; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2573 = io_dcache_ptw_pte_valid ? _GEN_2158 : _GEN_1498; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2574 = io_dcache_ptw_pte_valid ? _GEN_2159 : _GEN_1499; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2575 = io_dcache_ptw_pte_valid ? _GEN_2160 : _GEN_1500; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2576 = io_dcache_ptw_pte_valid ? _GEN_2161 : _GEN_1501; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2577 = io_dcache_ptw_pte_valid ? _GEN_2162 : _GEN_1502; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2578 = io_dcache_ptw_pte_valid ? _GEN_2163 : _GEN_1503; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2579 = io_dcache_ptw_pte_valid ? _GEN_2164 : _GEN_1504; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2580 = io_dcache_ptw_pte_valid ? _GEN_2165 : _GEN_1505; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2581 = io_dcache_ptw_pte_valid ? _GEN_2166 : _GEN_1506; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2582 = io_dcache_ptw_pte_valid ? _GEN_2167 : _GEN_1507; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2583 = io_dcache_ptw_pte_valid ? _GEN_2168 : _GEN_1508; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2584 = io_dcache_ptw_pte_valid ? _GEN_2169 : _GEN_1509; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2585 = io_dcache_ptw_pte_valid ? _GEN_2170 : _GEN_1510; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2586 = io_dcache_ptw_pte_valid ? _GEN_2171 : _GEN_1511; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2587 = io_dcache_ptw_pte_valid ? _GEN_2172 : _GEN_1512; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2588 = io_dcache_ptw_pte_valid ? _GEN_2173 : _GEN_1513; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2589 = io_dcache_ptw_pte_valid ? _GEN_2174 : _GEN_1514; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2590 = io_dcache_ptw_pte_valid ? _GEN_2175 : _GEN_1515; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2591 = io_dcache_ptw_pte_valid ? _GEN_2176 : _GEN_1516; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2592 = io_dcache_ptw_pte_valid ? _GEN_2177 : _GEN_1517; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2593 = io_dcache_ptw_pte_valid ? _GEN_2178 : _GEN_1518; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2594 = io_dcache_ptw_pte_valid ? _GEN_2179 : _GEN_1519; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2595 = io_dcache_ptw_pte_valid ? _GEN_2180 : _GEN_1520; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2596 = io_dcache_ptw_pte_valid ? _GEN_2181 : _GEN_1521; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2597 = io_dcache_ptw_pte_valid ? _GEN_2182 : _GEN_1522; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [15:0] _GEN_2598 = io_dcache_ptw_pte_valid ? _GEN_2183 : _GEN_1523; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2599 = io_dcache_ptw_pte_valid ? _GEN_2184 : _GEN_1524; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2600 = io_dcache_ptw_pte_valid ? _GEN_2185 : _GEN_1525; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2601 = io_dcache_ptw_pte_valid ? _GEN_2186 : _GEN_1526; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2602 = io_dcache_ptw_pte_valid ? _GEN_2187 : _GEN_1527; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2603 = io_dcache_ptw_pte_valid ? _GEN_2188 : _GEN_1528; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2604 = io_dcache_ptw_pte_valid ? _GEN_2189 : _GEN_1529; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2605 = io_dcache_ptw_pte_valid ? _GEN_2190 : _GEN_1530; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2606 = io_dcache_ptw_pte_valid ? _GEN_2191 : _GEN_1531; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2607 = io_dcache_ptw_pte_valid ? _GEN_2192 : _GEN_1532; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2608 = io_dcache_ptw_pte_valid ? _GEN_2193 : _GEN_1533; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2609 = io_dcache_ptw_pte_valid ? _GEN_2194 : _GEN_1534; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2610 = io_dcache_ptw_pte_valid ? _GEN_2195 : _GEN_1535; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2611 = io_dcache_ptw_pte_valid ? _GEN_2196 : _GEN_1536; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2612 = io_dcache_ptw_pte_valid ? _GEN_2197 : _GEN_1537; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2613 = io_dcache_ptw_pte_valid ? _GEN_2198 : _GEN_1538; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2614 = io_dcache_ptw_pte_valid ? _GEN_2199 : _GEN_1539; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2631 = io_dcache_ptw_pte_valid ? _GEN_2216 : _GEN_1556; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2632 = io_dcache_ptw_pte_valid ? _GEN_2217 : _GEN_1557; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2633 = io_dcache_ptw_pte_valid ? _GEN_2218 : _GEN_1558; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2634 = io_dcache_ptw_pte_valid ? _GEN_2219 : _GEN_1559; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2635 = io_dcache_ptw_pte_valid ? _GEN_2220 : _GEN_1560; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2636 = io_dcache_ptw_pte_valid ? _GEN_2221 : _GEN_1561; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2637 = io_dcache_ptw_pte_valid ? _GEN_2222 : _GEN_1562; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2638 = io_dcache_ptw_pte_valid ? _GEN_2223 : _GEN_1563; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2639 = io_dcache_ptw_pte_valid ? _GEN_2224 : _GEN_1564; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2640 = io_dcache_ptw_pte_valid ? _GEN_2225 : _GEN_1565; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2641 = io_dcache_ptw_pte_valid ? _GEN_2226 : _GEN_1566; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2642 = io_dcache_ptw_pte_valid ? _GEN_2227 : _GEN_1567; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2643 = io_dcache_ptw_pte_valid ? _GEN_2228 : _GEN_1568; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2644 = io_dcache_ptw_pte_valid ? _GEN_2229 : _GEN_1569; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2645 = io_dcache_ptw_pte_valid ? _GEN_2230 : _GEN_1570; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2646 = io_dcache_ptw_pte_valid ? _GEN_2231 : _GEN_1571; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2647 = io_dcache_ptw_pte_valid ? _GEN_2232 : _GEN_1572; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2648 = io_dcache_ptw_pte_valid ? _GEN_2233 : _GEN_1573; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2649 = io_dcache_ptw_pte_valid ? _GEN_2234 : _GEN_1574; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2650 = io_dcache_ptw_pte_valid ? _GEN_2235 : _GEN_1575; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2651 = io_dcache_ptw_pte_valid ? _GEN_2236 : _GEN_1576; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2652 = io_dcache_ptw_pte_valid ? _GEN_2237 : _GEN_1577; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2653 = io_dcache_ptw_pte_valid ? _GEN_2238 : _GEN_1578; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2654 = io_dcache_ptw_pte_valid ? _GEN_2239 : _GEN_1579; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2655 = io_dcache_ptw_pte_valid ? _GEN_2240 : _GEN_1580; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2656 = io_dcache_ptw_pte_valid ? _GEN_2241 : _GEN_1581; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2657 = io_dcache_ptw_pte_valid ? _GEN_2242 : _GEN_1582; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2658 = io_dcache_ptw_pte_valid ? _GEN_2243 : _GEN_1583; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2659 = io_dcache_ptw_pte_valid ? _GEN_2244 : _GEN_1584; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2660 = io_dcache_ptw_pte_valid ? _GEN_2245 : _GEN_1585; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2661 = io_dcache_ptw_pte_valid ? _GEN_2246 : _GEN_1586; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2662 = io_dcache_ptw_pte_valid ? _GEN_2247 : _GEN_1587; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2663 = io_dcache_ptw_pte_valid ? _GEN_2248 : _GEN_1588; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2664 = io_dcache_ptw_pte_valid ? _GEN_2249 : _GEN_1589; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2665 = io_dcache_ptw_pte_valid ? _GEN_2250 : _GEN_1590; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2666 = io_dcache_ptw_pte_valid ? _GEN_2251 : _GEN_1591; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2667 = io_dcache_ptw_pte_valid ? _GEN_2252 : _GEN_1592; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2668 = io_dcache_ptw_pte_valid ? _GEN_2253 : _GEN_1593; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2669 = io_dcache_ptw_pte_valid ? _GEN_2254 : _GEN_1594; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2670 = io_dcache_ptw_pte_valid ? _GEN_2255 : _GEN_1595; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2671 = io_dcache_ptw_pte_valid ? _GEN_2256 : _GEN_1596; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2672 = io_dcache_ptw_pte_valid ? _GEN_2257 : _GEN_1597; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2673 = io_dcache_ptw_pte_valid ? _GEN_2258 : _GEN_1598; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2674 = io_dcache_ptw_pte_valid ? _GEN_2259 : _GEN_1599; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2675 = io_dcache_ptw_pte_valid ? _GEN_2260 : _GEN_1600; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2676 = io_dcache_ptw_pte_valid ? _GEN_2261 : _GEN_1601; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2677 = io_dcache_ptw_pte_valid ? _GEN_2262 : _GEN_1602; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2678 = io_dcache_ptw_pte_valid ? _GEN_2263 : _GEN_1603; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2679 = io_dcache_ptw_pte_valid ? _GEN_2264 : _GEN_1604; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2680 = io_dcache_ptw_pte_valid ? _GEN_2265 : _GEN_1605; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2681 = io_dcache_ptw_pte_valid ? _GEN_2266 : _GEN_1606; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2682 = io_dcache_ptw_pte_valid ? _GEN_2267 : _GEN_1607; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2683 = io_dcache_ptw_pte_valid ? _GEN_2268 : _GEN_1608; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2684 = io_dcache_ptw_pte_valid ? _GEN_2269 : _GEN_1609; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2685 = io_dcache_ptw_pte_valid ? _GEN_2270 : _GEN_1610; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2686 = io_dcache_ptw_pte_valid ? _GEN_2271 : _GEN_1611; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2687 = io_dcache_ptw_pte_valid ? _GEN_2272 : _GEN_1612; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2688 = io_dcache_ptw_pte_valid ? _GEN_2273 : _GEN_1613; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2689 = io_dcache_ptw_pte_valid ? _GEN_2274 : _GEN_1614; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2690 = io_dcache_ptw_pte_valid ? _GEN_2275 : _GEN_1615; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2691 = io_dcache_ptw_pte_valid ? _GEN_2276 : _GEN_1616; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2692 = io_dcache_ptw_pte_valid ? _GEN_2277 : _GEN_1617; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2693 = io_dcache_ptw_pte_valid ? _GEN_2278 : _GEN_1618; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2694 = io_dcache_ptw_pte_valid ? _GEN_2279 : _GEN_1619; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2695 = io_dcache_ptw_pte_valid ? _GEN_2280 : _GEN_1620; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2696 = io_dcache_ptw_pte_valid ? _GEN_2281 : _GEN_1621; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2697 = io_dcache_ptw_pte_valid ? _GEN_2282 : _GEN_1622; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2698 = io_dcache_ptw_pte_valid ? _GEN_2283 : _GEN_1623; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2699 = io_dcache_ptw_pte_valid ? _GEN_2284 : _GEN_1624; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2700 = io_dcache_ptw_pte_valid ? _GEN_2285 : _GEN_1625; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2701 = io_dcache_ptw_pte_valid ? _GEN_2286 : _GEN_1626; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2702 = io_dcache_ptw_pte_valid ? _GEN_2287 : _GEN_1627; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2703 = io_dcache_ptw_pte_valid ? _GEN_2288 : _GEN_1628; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2704 = io_dcache_ptw_pte_valid ? _GEN_2289 : _GEN_1629; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2705 = io_dcache_ptw_pte_valid ? _GEN_2290 : _GEN_1630; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2706 = io_dcache_ptw_pte_valid ? _GEN_2291 : _GEN_1631; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2707 = io_dcache_ptw_pte_valid ? _GEN_2292 : _GEN_1632; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2708 = io_dcache_ptw_pte_valid ? _GEN_2293 : _GEN_1633; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2709 = io_dcache_ptw_pte_valid ? _GEN_2294 : _GEN_1634; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2710 = io_dcache_ptw_pte_valid ? _GEN_2295 : _GEN_1635; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2711 = io_dcache_ptw_pte_valid ? _GEN_2296 : _GEN_1636; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2712 = io_dcache_ptw_pte_valid ? _GEN_2297 : _GEN_1637; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2713 = io_dcache_ptw_pte_valid ? _GEN_2298 : _GEN_1638; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2714 = io_dcache_ptw_pte_valid ? _GEN_2299 : _GEN_1639; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2715 = io_dcache_ptw_pte_valid ? _GEN_2300 : _GEN_1640; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2716 = io_dcache_ptw_pte_valid ? _GEN_2301 : _GEN_1641; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2717 = io_dcache_ptw_pte_valid ? _GEN_2302 : _GEN_1642; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2718 = io_dcache_ptw_pte_valid ? _GEN_2303 : _GEN_1643; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2719 = io_dcache_ptw_pte_valid ? _GEN_2304 : _GEN_1644; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2720 = io_dcache_ptw_pte_valid ? _GEN_2305 : _GEN_1645; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2721 = io_dcache_ptw_pte_valid ? _GEN_2306 : _GEN_1646; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2722 = io_dcache_ptw_pte_valid ? _GEN_2307 : _GEN_1647; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2723 = io_dcache_ptw_pte_valid ? _GEN_2308 : _GEN_1648; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2724 = io_dcache_ptw_pte_valid ? _GEN_2309 : _GEN_1649; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2725 = io_dcache_ptw_pte_valid ? _GEN_2310 : _GEN_1650; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2726 = io_dcache_ptw_pte_valid ? _GEN_2311 : _GEN_1651; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2727 = io_dcache_ptw_pte_valid ? _GEN_2312 : _GEN_1652; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2728 = io_dcache_ptw_pte_valid ? _GEN_2313 : _GEN_1653; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2729 = io_dcache_ptw_pte_valid ? _GEN_2314 : _GEN_1654; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2730 = io_dcache_ptw_pte_valid ? _GEN_2315 : _GEN_1655; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2731 = io_dcache_ptw_pte_valid ? _GEN_2316 : _GEN_1656; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2732 = io_dcache_ptw_pte_valid ? _GEN_2317 : _GEN_1657; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2733 = io_dcache_ptw_pte_valid ? _GEN_2318 : _GEN_1658; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2734 = io_dcache_ptw_pte_valid ? _GEN_2319 : _GEN_1659; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2735 = io_dcache_ptw_pte_valid ? _GEN_2320 : _GEN_1660; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2736 = io_dcache_ptw_pte_valid ? _GEN_2321 : _GEN_1661; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2737 = io_dcache_ptw_pte_valid ? _GEN_2322 : _GEN_1662; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2738 = io_dcache_ptw_pte_valid ? _GEN_2323 : _GEN_1663; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2739 = io_dcache_ptw_pte_valid ? _GEN_2324 : _GEN_1664; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2740 = io_dcache_ptw_pte_valid ? _GEN_2325 : _GEN_1665; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2741 = io_dcache_ptw_pte_valid ? _GEN_2326 : _GEN_1666; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [19:0] _GEN_2742 = io_dcache_ptw_pte_valid ? _GEN_2327 : _GEN_1667; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2743 = io_dcache_ptw_pte_valid ? _GEN_2328 : _GEN_1668; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2744 = io_dcache_ptw_pte_valid ? _GEN_2329 : _GEN_1669; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2745 = io_dcache_ptw_pte_valid ? _GEN_2330 : _GEN_1670; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2746 = io_dcache_ptw_pte_valid ? _GEN_2331 : _GEN_1671; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2747 = io_dcache_ptw_pte_valid ? _GEN_2332 : _GEN_1672; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2748 = io_dcache_ptw_pte_valid ? _GEN_2333 : _GEN_1673; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2749 = io_dcache_ptw_pte_valid ? _GEN_2334 : _GEN_1674; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2750 = io_dcache_ptw_pte_valid ? _GEN_2335 : _GEN_1675; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2751 = io_dcache_ptw_pte_valid ? _GEN_2336 : _GEN_1676; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2752 = io_dcache_ptw_pte_valid ? _GEN_2337 : _GEN_1677; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2753 = io_dcache_ptw_pte_valid ? _GEN_2338 : _GEN_1678; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2754 = io_dcache_ptw_pte_valid ? _GEN_2339 : _GEN_1679; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2755 = io_dcache_ptw_pte_valid ? _GEN_2340 : _GEN_1680; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2756 = io_dcache_ptw_pte_valid ? _GEN_2341 : _GEN_1681; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2757 = io_dcache_ptw_pte_valid ? _GEN_2342 : _GEN_1682; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [17:0] _GEN_2758 = io_dcache_ptw_pte_valid ? _GEN_2343 : _GEN_1683; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire [26:0] _GEN_2759 = io_dcache_ptw_pte_valid ? _GEN_2344 : dtlb_vpn; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire [15:0] _GEN_2760 = io_dcache_ptw_pte_valid ? _GEN_2345 : dtlb_asid; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2761 = io_dcache_ptw_pte_valid ? _GEN_2346 : dtlb_flag_d; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2763 = io_dcache_ptw_pte_valid ? _GEN_2348 : dtlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2764 = io_dcache_ptw_pte_valid ? _GEN_2349 : dtlb_flag_u; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2765 = io_dcache_ptw_pte_valid ? _GEN_2350 : dtlb_flag_x; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2766 = io_dcache_ptw_pte_valid ? _GEN_2351 : dtlb_flag_w; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2767 = io_dcache_ptw_pte_valid ? _GEN_2352 : dtlb_flag_r; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire  _GEN_2768 = io_dcache_ptw_pte_valid ? _GEN_2353 : dtlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire [19:0] _GEN_2769 = io_dcache_ptw_pte_valid ? _GEN_2354 : dtlb_ppn; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire [17:0] _GEN_2770 = io_dcache_ptw_pte_valid ? _GEN_2355 : dtlb_rmask; // @[playground/src/cache/mmu/Tlb.scala 332:37 76:22]
  wire [3:0] _GEN_2771 = io_dcache_ptw_pte_valid ? _GEN_2356 : _GEN_1684; // @[playground/src/cache/mmu/Tlb.scala 332:37]
  wire  _GEN_2772 = io_dcache_complete_single_request ? 1'h0 : dpage_fault; // @[playground/src/cache/mmu/Tlb.scala 355:47 356:23 113:30]
  wire [1:0] _GEN_2774 = io_dcache_complete_single_request ? 2'h0 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 355:47 358:23 107:76]
  wire  _GEN_2775 = 2'h3 == dmmu_state ? _GEN_2772 : dpage_fault; // @[playground/src/cache/mmu/Tlb.scala 266:22 113:30]
  wire [1:0] _GEN_2777 = 2'h3 == dmmu_state ? _GEN_2774 : dmmu_state; // @[playground/src/cache/mmu/Tlb.scala 266:22 107:76]
  wire  _GEN_2926 = 2'h2 == dmmu_state ? _GEN_2711 : _GEN_1636; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2927 = 2'h2 == dmmu_state ? _GEN_2712 : _GEN_1637; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2928 = 2'h2 == dmmu_state ? _GEN_2713 : _GEN_1638; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2929 = 2'h2 == dmmu_state ? _GEN_2714 : _GEN_1639; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2930 = 2'h2 == dmmu_state ? _GEN_2715 : _GEN_1640; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2931 = 2'h2 == dmmu_state ? _GEN_2716 : _GEN_1641; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2932 = 2'h2 == dmmu_state ? _GEN_2717 : _GEN_1642; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2933 = 2'h2 == dmmu_state ? _GEN_2718 : _GEN_1643; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2934 = 2'h2 == dmmu_state ? _GEN_2719 : _GEN_1644; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2935 = 2'h2 == dmmu_state ? _GEN_2720 : _GEN_1645; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2936 = 2'h2 == dmmu_state ? _GEN_2721 : _GEN_1646; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2937 = 2'h2 == dmmu_state ? _GEN_2722 : _GEN_1647; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2938 = 2'h2 == dmmu_state ? _GEN_2723 : _GEN_1648; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2939 = 2'h2 == dmmu_state ? _GEN_2724 : _GEN_1649; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2940 = 2'h2 == dmmu_state ? _GEN_2725 : _GEN_1650; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2941 = 2'h2 == dmmu_state ? _GEN_2726 : _GEN_1651; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_2983 = 2'h2 == dmmu_state ? _GEN_2768 : dtlb_flag_v; // @[playground/src/cache/mmu/Tlb.scala 266:22 76:22]
  wire  _GEN_2997 = 2'h1 == dmmu_state ? _GEN_1955 : _GEN_2983; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3147 = 2'h1 == dmmu_state ? _GEN_1636 : _GEN_2926; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3148 = 2'h1 == dmmu_state ? _GEN_1637 : _GEN_2927; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3149 = 2'h1 == dmmu_state ? _GEN_1638 : _GEN_2928; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3150 = 2'h1 == dmmu_state ? _GEN_1639 : _GEN_2929; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3151 = 2'h1 == dmmu_state ? _GEN_1640 : _GEN_2930; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3152 = 2'h1 == dmmu_state ? _GEN_1641 : _GEN_2931; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3153 = 2'h1 == dmmu_state ? _GEN_1642 : _GEN_2932; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3154 = 2'h1 == dmmu_state ? _GEN_1643 : _GEN_2933; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3155 = 2'h1 == dmmu_state ? _GEN_1644 : _GEN_2934; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3156 = 2'h1 == dmmu_state ? _GEN_1645 : _GEN_2935; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3157 = 2'h1 == dmmu_state ? _GEN_1646 : _GEN_2936; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3158 = 2'h1 == dmmu_state ? _GEN_1647 : _GEN_2937; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3159 = 2'h1 == dmmu_state ? _GEN_1648 : _GEN_2938; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3160 = 2'h1 == dmmu_state ? _GEN_1649 : _GEN_2939; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3161 = 2'h1 == dmmu_state ? _GEN_1650 : _GEN_2940; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3162 = 2'h1 == dmmu_state ? _GEN_1651 : _GEN_2941; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3209 = 2'h0 == dmmu_state ? dtlb_flag_v : _GEN_2997; // @[playground/src/cache/mmu/Tlb.scala 266:22 76:22]
  wire  _GEN_3357 = 2'h0 == dmmu_state ? _GEN_1636 : _GEN_3147; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3358 = 2'h0 == dmmu_state ? _GEN_1637 : _GEN_3148; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3359 = 2'h0 == dmmu_state ? _GEN_1638 : _GEN_3149; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3360 = 2'h0 == dmmu_state ? _GEN_1639 : _GEN_3150; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3361 = 2'h0 == dmmu_state ? _GEN_1640 : _GEN_3151; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3362 = 2'h0 == dmmu_state ? _GEN_1641 : _GEN_3152; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3363 = 2'h0 == dmmu_state ? _GEN_1642 : _GEN_3153; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3364 = 2'h0 == dmmu_state ? _GEN_1643 : _GEN_3154; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3365 = 2'h0 == dmmu_state ? _GEN_1644 : _GEN_3155; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3366 = 2'h0 == dmmu_state ? _GEN_1645 : _GEN_3156; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3367 = 2'h0 == dmmu_state ? _GEN_1646 : _GEN_3157; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3368 = 2'h0 == dmmu_state ? _GEN_1647 : _GEN_3158; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3369 = 2'h0 == dmmu_state ? _GEN_1648 : _GEN_3159; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3370 = 2'h0 == dmmu_state ? _GEN_1649 : _GEN_3160; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3371 = 2'h0 == dmmu_state ? _GEN_1650 : _GEN_3161; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire  _GEN_3372 = 2'h0 == dmmu_state ? _GEN_1651 : _GEN_3162; // @[playground/src/cache/mmu/Tlb.scala 266:22]
  wire [14:0] src1 = io_sfence_vma_src_info_src1_data[26:12]; // @[playground/src/cache/mmu/Tlb.scala 364:46]
  wire [15:0] src2 = io_sfence_vma_src_info_src2_data[15:0]; // @[playground/src/cache/mmu/Tlb.scala 366:46]
  wire  _T_46 = |src1; // @[playground/src/cache/mmu/Tlb.scala 368:16]
  wire  _T_47 = ~(|src1); // @[playground/src/cache/mmu/Tlb.scala 368:10]
  wire  _T_48 = |src2; // @[playground/src/cache/mmu/Tlb.scala 368:29]
  wire  _T_49 = ~(|src2); // @[playground/src/cache/mmu/Tlb.scala 368:23]
  wire  _T_55 = itlb_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 377:22]
  wire  _T_56 = ~itlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 377:34]
  wire  _GEN_3406 = itlb_asid == src2 & ~itlb_flag_g ? 1'h0 : _GEN_1488; // @[playground/src/cache/mmu/Tlb.scala 377:48 378:21]
  wire  _T_58 = dtlb_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 380:22]
  wire  _T_59 = ~dtlb_flag_g; // @[playground/src/cache/mmu/Tlb.scala 380:34]
  wire  _GEN_3407 = dtlb_asid == src2 & ~dtlb_flag_g ? 1'h0 : _GEN_3209; // @[playground/src/cache/mmu/Tlb.scala 380:48 381:21]
  wire  _T_61 = tlbl2_0_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_62 = ~tlbl2_0_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3408 = tlbl2_0_asid == src2 & ~tlbl2_0_flag_g ? 1'h0 : _GEN_3357; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_64 = tlbl2_1_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_65 = ~tlbl2_1_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3409 = tlbl2_1_asid == src2 & ~tlbl2_1_flag_g ? 1'h0 : _GEN_3358; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_67 = tlbl2_2_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_68 = ~tlbl2_2_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3410 = tlbl2_2_asid == src2 & ~tlbl2_2_flag_g ? 1'h0 : _GEN_3359; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_70 = tlbl2_3_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_71 = ~tlbl2_3_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3411 = tlbl2_3_asid == src2 & ~tlbl2_3_flag_g ? 1'h0 : _GEN_3360; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_73 = tlbl2_4_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_74 = ~tlbl2_4_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3412 = tlbl2_4_asid == src2 & ~tlbl2_4_flag_g ? 1'h0 : _GEN_3361; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_76 = tlbl2_5_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_77 = ~tlbl2_5_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3413 = tlbl2_5_asid == src2 & ~tlbl2_5_flag_g ? 1'h0 : _GEN_3362; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_79 = tlbl2_6_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_80 = ~tlbl2_6_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3414 = tlbl2_6_asid == src2 & ~tlbl2_6_flag_g ? 1'h0 : _GEN_3363; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_82 = tlbl2_7_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_83 = ~tlbl2_7_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3415 = tlbl2_7_asid == src2 & ~tlbl2_7_flag_g ? 1'h0 : _GEN_3364; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_85 = tlbl2_8_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_86 = ~tlbl2_8_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3416 = tlbl2_8_asid == src2 & ~tlbl2_8_flag_g ? 1'h0 : _GEN_3365; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_88 = tlbl2_9_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_89 = ~tlbl2_9_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3417 = tlbl2_9_asid == src2 & ~tlbl2_9_flag_g ? 1'h0 : _GEN_3366; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_91 = tlbl2_10_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_92 = ~tlbl2_10_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3418 = tlbl2_10_asid == src2 & ~tlbl2_10_flag_g ? 1'h0 : _GEN_3367; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_94 = tlbl2_11_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_95 = ~tlbl2_11_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3419 = tlbl2_11_asid == src2 & ~tlbl2_11_flag_g ? 1'h0 : _GEN_3368; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_97 = tlbl2_12_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_98 = ~tlbl2_12_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3420 = tlbl2_12_asid == src2 & ~tlbl2_12_flag_g ? 1'h0 : _GEN_3369; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_100 = tlbl2_13_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_101 = ~tlbl2_13_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3421 = tlbl2_13_asid == src2 & ~tlbl2_13_flag_g ? 1'h0 : _GEN_3370; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_103 = tlbl2_14_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_104 = ~tlbl2_14_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3422 = tlbl2_14_asid == src2 & ~tlbl2_14_flag_g ? 1'h0 : _GEN_3371; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire  _T_106 = tlbl2_15_asid == src2; // @[playground/src/cache/mmu/Tlb.scala 384:28]
  wire  _T_107 = ~tlbl2_15_flag_g; // @[playground/src/cache/mmu/Tlb.scala 384:40]
  wire  _GEN_3423 = tlbl2_15_asid == src2 & ~tlbl2_15_flag_g ? 1'h0 : _GEN_3372; // @[playground/src/cache/mmu/Tlb.scala 384:58 385:27]
  wire [26:0] _GEN_3550 = {{12'd0}, src1}; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire [26:0] _T_113 = _GEN_3550 & itlbl1_hit_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_115 = _T_113 == _itlbl1_hit_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3424 = _T_115 ? 1'h0 : _GEN_1488; // @[playground/src/cache/mmu/Tlb.scala 390:47 391:21]
  wire [26:0] _T_116 = _GEN_3550 & dtlbl1_hit_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_118 = _T_116 == _dtlbl1_hit_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3425 = _T_118 ? 1'h0 : _GEN_3209; // @[playground/src/cache/mmu/Tlb.scala 393:47 394:21]
  wire [26:0] _T_119 = _GEN_3550 & il2_hit_vec_fullmask; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_121 = _T_119 == _il2_hit_vec_T_1; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3426 = _T_121 ? 1'h0 : _GEN_3357; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_122 = _GEN_3550 & il2_hit_vec_fullmask_1; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_124 = _T_122 == _il2_hit_vec_T_8; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3427 = _T_124 ? 1'h0 : _GEN_3358; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_125 = _GEN_3550 & il2_hit_vec_fullmask_2; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_127 = _T_125 == _il2_hit_vec_T_15; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3428 = _T_127 ? 1'h0 : _GEN_3359; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_128 = _GEN_3550 & il2_hit_vec_fullmask_3; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_130 = _T_128 == _il2_hit_vec_T_22; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3429 = _T_130 ? 1'h0 : _GEN_3360; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_131 = _GEN_3550 & il2_hit_vec_fullmask_4; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_133 = _T_131 == _il2_hit_vec_T_29; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3430 = _T_133 ? 1'h0 : _GEN_3361; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_134 = _GEN_3550 & il2_hit_vec_fullmask_5; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_136 = _T_134 == _il2_hit_vec_T_36; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3431 = _T_136 ? 1'h0 : _GEN_3362; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_137 = _GEN_3550 & il2_hit_vec_fullmask_6; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_139 = _T_137 == _il2_hit_vec_T_43; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3432 = _T_139 ? 1'h0 : _GEN_3363; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_140 = _GEN_3550 & il2_hit_vec_fullmask_7; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_142 = _T_140 == _il2_hit_vec_T_50; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3433 = _T_142 ? 1'h0 : _GEN_3364; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_143 = _GEN_3550 & il2_hit_vec_fullmask_8; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_145 = _T_143 == _il2_hit_vec_T_57; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3434 = _T_145 ? 1'h0 : _GEN_3365; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_146 = _GEN_3550 & il2_hit_vec_fullmask_9; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_148 = _T_146 == _il2_hit_vec_T_64; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3435 = _T_148 ? 1'h0 : _GEN_3366; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_149 = _GEN_3550 & il2_hit_vec_fullmask_10; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_151 = _T_149 == _il2_hit_vec_T_71; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3436 = _T_151 ? 1'h0 : _GEN_3367; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_152 = _GEN_3550 & il2_hit_vec_fullmask_11; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_154 = _T_152 == _il2_hit_vec_T_78; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3437 = _T_154 ? 1'h0 : _GEN_3368; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_155 = _GEN_3550 & il2_hit_vec_fullmask_12; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_157 = _T_155 == _il2_hit_vec_T_85; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3438 = _T_157 ? 1'h0 : _GEN_3369; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_158 = _GEN_3550 & il2_hit_vec_fullmask_13; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_160 = _T_158 == _il2_hit_vec_T_92; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3439 = _T_160 ? 1'h0 : _GEN_3370; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_161 = _GEN_3550 & il2_hit_vec_fullmask_14; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_163 = _T_161 == _il2_hit_vec_T_99; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3440 = _T_163 ? 1'h0 : _GEN_3371; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire [26:0] _T_164 = _GEN_3550 & il2_hit_vec_fullmask_15; // @[playground/src/defines/TlbBundles.scala 37:10]
  wire  _T_166 = _T_164 == _il2_hit_vec_T_106; // @[playground/src/defines/TlbBundles.scala 37:22]
  wire  _GEN_3441 = _T_166 ? 1'h0 : _GEN_3372; // @[playground/src/cache/mmu/Tlb.scala 397:57 398:27]
  wire  _GEN_3442 = _T_55 & _T_115 & _T_56 ? 1'h0 : _GEN_1488; // @[playground/src/cache/mmu/Tlb.scala 403:85 404:21]
  wire  _GEN_3443 = _T_58 & _T_118 & _T_59 ? 1'h0 : _GEN_3209; // @[playground/src/cache/mmu/Tlb.scala 406:85 407:21]
  wire  _GEN_3444 = _T_61 & _T_121 & _T_62 ? 1'h0 : _GEN_3357; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3445 = _T_64 & _T_124 & _T_65 ? 1'h0 : _GEN_3358; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3446 = _T_67 & _T_127 & _T_68 ? 1'h0 : _GEN_3359; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3447 = _T_70 & _T_130 & _T_71 ? 1'h0 : _GEN_3360; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3448 = _T_73 & _T_133 & _T_74 ? 1'h0 : _GEN_3361; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3449 = _T_76 & _T_136 & _T_77 ? 1'h0 : _GEN_3362; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3450 = _T_79 & _T_139 & _T_80 ? 1'h0 : _GEN_3363; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3451 = _T_82 & _T_142 & _T_83 ? 1'h0 : _GEN_3364; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3452 = _T_85 & _T_145 & _T_86 ? 1'h0 : _GEN_3365; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3453 = _T_88 & _T_148 & _T_89 ? 1'h0 : _GEN_3366; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3454 = _T_91 & _T_151 & _T_92 ? 1'h0 : _GEN_3367; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3455 = _T_94 & _T_154 & _T_95 ? 1'h0 : _GEN_3368; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3456 = _T_97 & _T_157 & _T_98 ? 1'h0 : _GEN_3369; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3457 = _T_100 & _T_160 & _T_101 ? 1'h0 : _GEN_3370; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3458 = _T_103 & _T_163 & _T_104 ? 1'h0 : _GEN_3371; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3459 = _T_106 & _T_166 & _T_107 ? 1'h0 : _GEN_3372; // @[playground/src/cache/mmu/Tlb.scala 410:103 411:27]
  wire  _GEN_3460 = _T_46 & _T_48 ? _GEN_3442 : _GEN_1488; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3461 = _T_46 & _T_48 ? _GEN_3443 : _GEN_3209; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3462 = _T_46 & _T_48 ? _GEN_3444 : _GEN_3357; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3463 = _T_46 & _T_48 ? _GEN_3445 : _GEN_3358; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3464 = _T_46 & _T_48 ? _GEN_3446 : _GEN_3359; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3465 = _T_46 & _T_48 ? _GEN_3447 : _GEN_3360; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3466 = _T_46 & _T_48 ? _GEN_3448 : _GEN_3361; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3467 = _T_46 & _T_48 ? _GEN_3449 : _GEN_3362; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3468 = _T_46 & _T_48 ? _GEN_3450 : _GEN_3363; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3469 = _T_46 & _T_48 ? _GEN_3451 : _GEN_3364; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3470 = _T_46 & _T_48 ? _GEN_3452 : _GEN_3365; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3471 = _T_46 & _T_48 ? _GEN_3453 : _GEN_3366; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3472 = _T_46 & _T_48 ? _GEN_3454 : _GEN_3367; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3473 = _T_46 & _T_48 ? _GEN_3455 : _GEN_3368; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3474 = _T_46 & _T_48 ? _GEN_3456 : _GEN_3369; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3475 = _T_46 & _T_48 ? _GEN_3457 : _GEN_3370; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3476 = _T_46 & _T_48 ? _GEN_3458 : _GEN_3371; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3477 = _T_46 & _T_48 ? _GEN_3459 : _GEN_3372; // @[playground/src/cache/mmu/Tlb.scala 401:38]
  wire  _GEN_3478 = _T_46 & _T_49 ? _GEN_3424 : _GEN_3460; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3479 = _T_46 & _T_49 ? _GEN_3425 : _GEN_3461; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3480 = _T_46 & _T_49 ? _GEN_3426 : _GEN_3462; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3481 = _T_46 & _T_49 ? _GEN_3427 : _GEN_3463; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3482 = _T_46 & _T_49 ? _GEN_3428 : _GEN_3464; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3483 = _T_46 & _T_49 ? _GEN_3429 : _GEN_3465; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3484 = _T_46 & _T_49 ? _GEN_3430 : _GEN_3466; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3485 = _T_46 & _T_49 ? _GEN_3431 : _GEN_3467; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3486 = _T_46 & _T_49 ? _GEN_3432 : _GEN_3468; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3487 = _T_46 & _T_49 ? _GEN_3433 : _GEN_3469; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3488 = _T_46 & _T_49 ? _GEN_3434 : _GEN_3470; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3489 = _T_46 & _T_49 ? _GEN_3435 : _GEN_3471; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3490 = _T_46 & _T_49 ? _GEN_3436 : _GEN_3472; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3491 = _T_46 & _T_49 ? _GEN_3437 : _GEN_3473; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3492 = _T_46 & _T_49 ? _GEN_3438 : _GEN_3474; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3493 = _T_46 & _T_49 ? _GEN_3439 : _GEN_3475; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3494 = _T_46 & _T_49 ? _GEN_3440 : _GEN_3476; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire  _GEN_3495 = _T_46 & _T_49 ? _GEN_3441 : _GEN_3477; // @[playground/src/cache/mmu/Tlb.scala 388:39]
  wire [19:0] imasktag_fullmask = {2'h3,itlb_rmask}; // @[playground/src/defines/TlbBundles.scala 41:23]
  wire [19:0] _imasktag_T = itlb_ppn & imasktag_fullmask; // @[playground/src/defines/TlbBundles.scala 42:10]
  wire [19:0] _imasktag_T_1 = ~imasktag_fullmask; // @[playground/src/defines/TlbBundles.scala 42:31]
  wire [26:0] _GEN_3586 = {{7'd0}, _imasktag_T_1}; // @[playground/src/defines/TlbBundles.scala 42:29]
  wire [26:0] _imasktag_T_2 = ivpn & _GEN_3586; // @[playground/src/defines/TlbBundles.scala 42:29]
  wire [26:0] _GEN_3587 = {{7'd0}, _imasktag_T}; // @[playground/src/defines/TlbBundles.scala 42:22]
  wire [26:0] imasktag = _GEN_3587 | _imasktag_T_2; // @[playground/src/defines/TlbBundles.scala 42:22]
  wire [19:0] dmasktag_fullmask = {2'h3,dtlb_rmask}; // @[playground/src/defines/TlbBundles.scala 41:23]
  wire [19:0] _dmasktag_T = dtlb_ppn & dmasktag_fullmask; // @[playground/src/defines/TlbBundles.scala 42:10]
  wire [19:0] _dmasktag_T_1 = ~dmasktag_fullmask; // @[playground/src/defines/TlbBundles.scala 42:31]
  wire [26:0] _GEN_3588 = {{7'd0}, _dmasktag_T_1}; // @[playground/src/defines/TlbBundles.scala 42:29]
  wire [26:0] _dmasktag_T_2 = dvpn & _GEN_3588; // @[playground/src/defines/TlbBundles.scala 42:29]
  wire [26:0] _GEN_3589 = {{7'd0}, _dmasktag_T}; // @[playground/src/defines/TlbBundles.scala 42:22]
  wire [26:0] dmasktag = _GEN_3589 | _dmasktag_T_2; // @[playground/src/defines/TlbBundles.scala 42:22]
  wire [63:0] _io_icache_uncached_T = io_icache_vaddr ^ 64'h30000000; // @[playground/src/defines/Const.scala 78:13]
  wire  _io_icache_uncached_T_2 = _io_icache_uncached_T[31:28] == 4'h0; // @[playground/src/defines/Const.scala 78:48]
  wire [63:0] _io_icache_uncached_T_3 = io_icache_vaddr ^ 64'h40000000; // @[playground/src/defines/Const.scala 78:13]
  wire  _io_icache_uncached_T_5 = _io_icache_uncached_T_3[31:30] == 2'h0; // @[playground/src/defines/Const.scala 78:48]
  wire [26:0] _io_icache_ptag_T = ivm_enabled ? imasktag : ivpn; // @[playground/src/cache/mmu/Tlb.scala 421:28]
  wire [63:0] _io_dcache_uncached_T = io_dcache_vaddr ^ 64'h30000000; // @[playground/src/defines/Const.scala 78:13]
  wire  _io_dcache_uncached_T_2 = _io_dcache_uncached_T[31:28] == 4'h0; // @[playground/src/defines/Const.scala 78:48]
  wire [63:0] _io_dcache_uncached_T_3 = io_dcache_vaddr ^ 64'h40000000; // @[playground/src/defines/Const.scala 78:13]
  wire  _io_dcache_uncached_T_5 = _io_dcache_uncached_T_3[31:30] == 2'h0; // @[playground/src/defines/Const.scala 78:48]
  wire [26:0] _io_dcache_ptag_T = dvm_enabled ? dmasktag : dvpn; // @[playground/src/cache/mmu/Tlb.scala 425:28]
  assign io_icache_uncached = _io_icache_uncached_T_2 | _io_icache_uncached_T_5; // @[playground/src/defines/Const.scala 80:15]
  assign io_icache_hit = 2'h0 == immu_state & _GEN_27; // @[playground/src/cache/mmu/Tlb.scala 193:22 134:26]
  assign io_icache_ptag = _io_icache_ptag_T[19:0]; // @[playground/src/cache/mmu/Tlb.scala 421:22]
  assign io_icache_paddr = {io_icache_ptag,io_icache_vaddr[11:0]}; // @[playground/src/cache/mmu/Tlb.scala 422:28]
  assign io_icache_page_fault = ipage_fault; // @[playground/src/cache/mmu/Tlb.scala 138:26]
  assign io_dcache_uncached = _io_dcache_uncached_T_2 | _io_dcache_uncached_T_5; // @[playground/src/defines/Const.scala 80:15]
  assign io_dcache_hit = 2'h0 == dmmu_state & _GEN_1750; // @[playground/src/cache/mmu/Tlb.scala 266:22 135:26]
  assign io_dcache_ptag = _io_dcache_ptag_T[19:0]; // @[playground/src/cache/mmu/Tlb.scala 425:22]
  assign io_dcache_paddr = {io_dcache_ptag,io_dcache_vaddr[11:0]}; // @[playground/src/cache/mmu/Tlb.scala 426:28]
  assign io_dcache_page_fault = dpage_fault; // @[playground/src/cache/mmu/Tlb.scala 139:26]
  assign io_dcache_ptw_vpn_valid = choose_icache ? req_ptw_0 : req_ptw_1; // @[playground/src/cache/mmu/Tlb.scala 142:35]
  assign io_dcache_ptw_vpn_bits = choose_icache ? ivpn : dvpn; // @[playground/src/cache/mmu/Tlb.scala 144:35]
  assign io_dcache_ptw_access_type = choose_icache ? 2'h0 : io_dcache_access_type; // @[playground/src/cache/mmu/Tlb.scala 143:35]
  assign io_dcache_csr_satp = io_csr_satp; // @[playground/src/cache/mmu/Tlb.scala 146:17]
  assign io_dcache_csr_mstatus = io_csr_mstatus; // @[playground/src/cache/mmu/Tlb.scala 146:17]
  assign io_dcache_csr_imode = io_csr_imode; // @[playground/src/cache/mmu/Tlb.scala 146:17]
  assign io_dcache_csr_dmode = io_csr_dmode; // @[playground/src/cache/mmu/Tlb.scala 146:17]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_vpn <= _GEN_44; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_vpn <= _GEN_1038;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_asid <= _GEN_60; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_asid <= _GEN_1039;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_flag_g <= _GEN_108; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_flag_g <= _GEN_1042;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_flag_u <= _GEN_124; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_flag_u <= _GEN_1043;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_flag_x <= _GEN_140; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_flag_x <= _GEN_1044;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        itlb_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 370:19]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        itlb_flag_v <= _GEN_3406;
      end else begin
        itlb_flag_v <= _GEN_3478;
      end
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_flag_v <= _GEN_232;
      end else begin
        itlb_flag_v <= _GEN_1262;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_ppn <= _GEN_204; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_ppn <= _GEN_1048;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 75:22]
      itlb_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 75:22]
    end else if (!(2'h0 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
          itlb_rmask <= _GEN_220; // @[playground/src/cache/mmu/Tlb.scala 222:20]
        end
      end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        itlb_rmask <= _GEN_1049;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_vpn <= _GEN_1767; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_vpn <= _GEN_2759;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_asid <= _GEN_1783; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_asid <= _GEN_2760;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_flag_d <= _GEN_1799; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_d <= _GEN_2761;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_flag_g <= _GEN_1831; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_g <= _GEN_2763;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_flag_u <= _GEN_1847; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_u <= _GEN_2764;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_flag_x <= _GEN_1863; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_x <= _GEN_2765;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_flag_w <= _GEN_1879; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_w <= _GEN_2766;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_flag_r <= _GEN_1895; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_r <= _GEN_2767;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        dtlb_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 371:19]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        dtlb_flag_v <= _GEN_3407;
      end else begin
        dtlb_flag_v <= _GEN_3479;
      end
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_flag_v <= _GEN_1955;
      end else begin
        dtlb_flag_v <= _GEN_2983;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_ppn <= _GEN_1927; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_ppn <= _GEN_2769;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 76:22]
      dtlb_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 76:22]
    end else if (!(2'h0 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
          dtlb_rmask <= _GEN_1943; // @[playground/src/cache/mmu/Tlb.scala 322:20]
        end
      end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dtlb_rmask <= _GEN_2770;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_vpn <= _GEN_1492;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_vpn <= _GEN_1492;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_vpn <= _GEN_2567;
    end else begin
      tlbl2_0_vpn <= _GEN_1492;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_asid <= _GEN_1508;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_asid <= _GEN_1508;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_asid <= _GEN_2583;
    end else begin
      tlbl2_0_asid <= _GEN_1508;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_d <= _GEN_1524;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_d <= _GEN_1524;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_d <= _GEN_2599;
    end else begin
      tlbl2_0_flag_d <= _GEN_1524;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_g <= _GEN_1556;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_g <= _GEN_1556;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_g <= _GEN_2631;
    end else begin
      tlbl2_0_flag_g <= _GEN_1556;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_u <= _GEN_1572;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_u <= _GEN_1572;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_u <= _GEN_2647;
    end else begin
      tlbl2_0_flag_u <= _GEN_1572;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_x <= _GEN_1588;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_x <= _GEN_1588;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_x <= _GEN_2663;
    end else begin
      tlbl2_0_flag_x <= _GEN_1588;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_w <= _GEN_1604;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_w <= _GEN_1604;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_w <= _GEN_2679;
    end else begin
      tlbl2_0_flag_w <= _GEN_1604;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_r <= _GEN_1620;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_r <= _GEN_1620;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_r <= _GEN_2695;
    end else begin
      tlbl2_0_flag_r <= _GEN_1620;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_0_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_0_flag_v <= _GEN_3408;
      end else begin
        tlbl2_0_flag_v <= _GEN_3480;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_v <= _GEN_1636;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_flag_v <= _GEN_1636;
    end else begin
      tlbl2_0_flag_v <= _GEN_2926;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_ppn <= _GEN_1652;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_ppn <= _GEN_1652;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_ppn <= _GEN_2727;
    end else begin
      tlbl2_0_ppn <= _GEN_1652;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_0_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_rmask <= _GEN_1668;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_rmask <= _GEN_1668;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_0_rmask <= _GEN_2743;
    end else begin
      tlbl2_0_rmask <= _GEN_1668;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_vpn <= _GEN_1493;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_vpn <= _GEN_1493;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_vpn <= _GEN_2568;
    end else begin
      tlbl2_1_vpn <= _GEN_1493;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_asid <= _GEN_1509;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_asid <= _GEN_1509;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_asid <= _GEN_2584;
    end else begin
      tlbl2_1_asid <= _GEN_1509;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_d <= _GEN_1525;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_d <= _GEN_1525;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_d <= _GEN_2600;
    end else begin
      tlbl2_1_flag_d <= _GEN_1525;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_g <= _GEN_1557;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_g <= _GEN_1557;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_g <= _GEN_2632;
    end else begin
      tlbl2_1_flag_g <= _GEN_1557;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_u <= _GEN_1573;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_u <= _GEN_1573;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_u <= _GEN_2648;
    end else begin
      tlbl2_1_flag_u <= _GEN_1573;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_x <= _GEN_1589;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_x <= _GEN_1589;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_x <= _GEN_2664;
    end else begin
      tlbl2_1_flag_x <= _GEN_1589;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_w <= _GEN_1605;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_w <= _GEN_1605;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_w <= _GEN_2680;
    end else begin
      tlbl2_1_flag_w <= _GEN_1605;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_r <= _GEN_1621;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_r <= _GEN_1621;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_r <= _GEN_2696;
    end else begin
      tlbl2_1_flag_r <= _GEN_1621;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_1_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_1_flag_v <= _GEN_3409;
      end else begin
        tlbl2_1_flag_v <= _GEN_3481;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_v <= _GEN_1637;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_flag_v <= _GEN_1637;
    end else begin
      tlbl2_1_flag_v <= _GEN_2927;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_ppn <= _GEN_1653;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_ppn <= _GEN_1653;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_ppn <= _GEN_2728;
    end else begin
      tlbl2_1_ppn <= _GEN_1653;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_1_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_rmask <= _GEN_1669;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_rmask <= _GEN_1669;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_1_rmask <= _GEN_2744;
    end else begin
      tlbl2_1_rmask <= _GEN_1669;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_vpn <= _GEN_1494;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_vpn <= _GEN_1494;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_vpn <= _GEN_2569;
    end else begin
      tlbl2_2_vpn <= _GEN_1494;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_asid <= _GEN_1510;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_asid <= _GEN_1510;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_asid <= _GEN_2585;
    end else begin
      tlbl2_2_asid <= _GEN_1510;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_d <= _GEN_1526;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_d <= _GEN_1526;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_d <= _GEN_2601;
    end else begin
      tlbl2_2_flag_d <= _GEN_1526;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_g <= _GEN_1558;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_g <= _GEN_1558;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_g <= _GEN_2633;
    end else begin
      tlbl2_2_flag_g <= _GEN_1558;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_u <= _GEN_1574;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_u <= _GEN_1574;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_u <= _GEN_2649;
    end else begin
      tlbl2_2_flag_u <= _GEN_1574;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_x <= _GEN_1590;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_x <= _GEN_1590;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_x <= _GEN_2665;
    end else begin
      tlbl2_2_flag_x <= _GEN_1590;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_w <= _GEN_1606;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_w <= _GEN_1606;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_w <= _GEN_2681;
    end else begin
      tlbl2_2_flag_w <= _GEN_1606;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_r <= _GEN_1622;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_r <= _GEN_1622;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_r <= _GEN_2697;
    end else begin
      tlbl2_2_flag_r <= _GEN_1622;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_2_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_2_flag_v <= _GEN_3410;
      end else begin
        tlbl2_2_flag_v <= _GEN_3482;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_v <= _GEN_1638;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_flag_v <= _GEN_1638;
    end else begin
      tlbl2_2_flag_v <= _GEN_2928;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_ppn <= _GEN_1654;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_ppn <= _GEN_1654;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_ppn <= _GEN_2729;
    end else begin
      tlbl2_2_ppn <= _GEN_1654;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_2_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_rmask <= _GEN_1670;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_rmask <= _GEN_1670;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_2_rmask <= _GEN_2745;
    end else begin
      tlbl2_2_rmask <= _GEN_1670;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_vpn <= _GEN_1495;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_vpn <= _GEN_1495;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_vpn <= _GEN_2570;
    end else begin
      tlbl2_3_vpn <= _GEN_1495;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_asid <= _GEN_1511;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_asid <= _GEN_1511;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_asid <= _GEN_2586;
    end else begin
      tlbl2_3_asid <= _GEN_1511;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_d <= _GEN_1527;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_d <= _GEN_1527;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_d <= _GEN_2602;
    end else begin
      tlbl2_3_flag_d <= _GEN_1527;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_g <= _GEN_1559;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_g <= _GEN_1559;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_g <= _GEN_2634;
    end else begin
      tlbl2_3_flag_g <= _GEN_1559;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_u <= _GEN_1575;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_u <= _GEN_1575;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_u <= _GEN_2650;
    end else begin
      tlbl2_3_flag_u <= _GEN_1575;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_x <= _GEN_1591;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_x <= _GEN_1591;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_x <= _GEN_2666;
    end else begin
      tlbl2_3_flag_x <= _GEN_1591;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_w <= _GEN_1607;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_w <= _GEN_1607;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_w <= _GEN_2682;
    end else begin
      tlbl2_3_flag_w <= _GEN_1607;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_r <= _GEN_1623;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_r <= _GEN_1623;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_r <= _GEN_2698;
    end else begin
      tlbl2_3_flag_r <= _GEN_1623;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_3_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_3_flag_v <= _GEN_3411;
      end else begin
        tlbl2_3_flag_v <= _GEN_3483;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_v <= _GEN_1639;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_flag_v <= _GEN_1639;
    end else begin
      tlbl2_3_flag_v <= _GEN_2929;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_ppn <= _GEN_1655;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_ppn <= _GEN_1655;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_ppn <= _GEN_2730;
    end else begin
      tlbl2_3_ppn <= _GEN_1655;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_3_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_rmask <= _GEN_1671;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_rmask <= _GEN_1671;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_3_rmask <= _GEN_2746;
    end else begin
      tlbl2_3_rmask <= _GEN_1671;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_vpn <= _GEN_1496;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_vpn <= _GEN_1496;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_vpn <= _GEN_2571;
    end else begin
      tlbl2_4_vpn <= _GEN_1496;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_asid <= _GEN_1512;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_asid <= _GEN_1512;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_asid <= _GEN_2587;
    end else begin
      tlbl2_4_asid <= _GEN_1512;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_d <= _GEN_1528;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_d <= _GEN_1528;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_d <= _GEN_2603;
    end else begin
      tlbl2_4_flag_d <= _GEN_1528;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_g <= _GEN_1560;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_g <= _GEN_1560;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_g <= _GEN_2635;
    end else begin
      tlbl2_4_flag_g <= _GEN_1560;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_u <= _GEN_1576;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_u <= _GEN_1576;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_u <= _GEN_2651;
    end else begin
      tlbl2_4_flag_u <= _GEN_1576;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_x <= _GEN_1592;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_x <= _GEN_1592;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_x <= _GEN_2667;
    end else begin
      tlbl2_4_flag_x <= _GEN_1592;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_w <= _GEN_1608;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_w <= _GEN_1608;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_w <= _GEN_2683;
    end else begin
      tlbl2_4_flag_w <= _GEN_1608;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_r <= _GEN_1624;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_r <= _GEN_1624;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_r <= _GEN_2699;
    end else begin
      tlbl2_4_flag_r <= _GEN_1624;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_4_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_4_flag_v <= _GEN_3412;
      end else begin
        tlbl2_4_flag_v <= _GEN_3484;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_v <= _GEN_1640;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_flag_v <= _GEN_1640;
    end else begin
      tlbl2_4_flag_v <= _GEN_2930;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_ppn <= _GEN_1656;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_ppn <= _GEN_1656;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_ppn <= _GEN_2731;
    end else begin
      tlbl2_4_ppn <= _GEN_1656;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_4_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_rmask <= _GEN_1672;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_rmask <= _GEN_1672;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_4_rmask <= _GEN_2747;
    end else begin
      tlbl2_4_rmask <= _GEN_1672;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_vpn <= _GEN_1497;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_vpn <= _GEN_1497;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_vpn <= _GEN_2572;
    end else begin
      tlbl2_5_vpn <= _GEN_1497;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_asid <= _GEN_1513;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_asid <= _GEN_1513;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_asid <= _GEN_2588;
    end else begin
      tlbl2_5_asid <= _GEN_1513;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_d <= _GEN_1529;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_d <= _GEN_1529;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_d <= _GEN_2604;
    end else begin
      tlbl2_5_flag_d <= _GEN_1529;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_g <= _GEN_1561;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_g <= _GEN_1561;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_g <= _GEN_2636;
    end else begin
      tlbl2_5_flag_g <= _GEN_1561;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_u <= _GEN_1577;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_u <= _GEN_1577;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_u <= _GEN_2652;
    end else begin
      tlbl2_5_flag_u <= _GEN_1577;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_x <= _GEN_1593;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_x <= _GEN_1593;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_x <= _GEN_2668;
    end else begin
      tlbl2_5_flag_x <= _GEN_1593;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_w <= _GEN_1609;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_w <= _GEN_1609;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_w <= _GEN_2684;
    end else begin
      tlbl2_5_flag_w <= _GEN_1609;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_r <= _GEN_1625;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_r <= _GEN_1625;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_r <= _GEN_2700;
    end else begin
      tlbl2_5_flag_r <= _GEN_1625;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_5_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_5_flag_v <= _GEN_3413;
      end else begin
        tlbl2_5_flag_v <= _GEN_3485;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_v <= _GEN_1641;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_flag_v <= _GEN_1641;
    end else begin
      tlbl2_5_flag_v <= _GEN_2931;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_ppn <= _GEN_1657;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_ppn <= _GEN_1657;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_ppn <= _GEN_2732;
    end else begin
      tlbl2_5_ppn <= _GEN_1657;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_5_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_rmask <= _GEN_1673;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_rmask <= _GEN_1673;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_5_rmask <= _GEN_2748;
    end else begin
      tlbl2_5_rmask <= _GEN_1673;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_vpn <= _GEN_1498;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_vpn <= _GEN_1498;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_vpn <= _GEN_2573;
    end else begin
      tlbl2_6_vpn <= _GEN_1498;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_asid <= _GEN_1514;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_asid <= _GEN_1514;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_asid <= _GEN_2589;
    end else begin
      tlbl2_6_asid <= _GEN_1514;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_d <= _GEN_1530;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_d <= _GEN_1530;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_d <= _GEN_2605;
    end else begin
      tlbl2_6_flag_d <= _GEN_1530;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_g <= _GEN_1562;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_g <= _GEN_1562;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_g <= _GEN_2637;
    end else begin
      tlbl2_6_flag_g <= _GEN_1562;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_u <= _GEN_1578;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_u <= _GEN_1578;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_u <= _GEN_2653;
    end else begin
      tlbl2_6_flag_u <= _GEN_1578;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_x <= _GEN_1594;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_x <= _GEN_1594;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_x <= _GEN_2669;
    end else begin
      tlbl2_6_flag_x <= _GEN_1594;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_w <= _GEN_1610;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_w <= _GEN_1610;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_w <= _GEN_2685;
    end else begin
      tlbl2_6_flag_w <= _GEN_1610;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_r <= _GEN_1626;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_r <= _GEN_1626;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_r <= _GEN_2701;
    end else begin
      tlbl2_6_flag_r <= _GEN_1626;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_6_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_6_flag_v <= _GEN_3414;
      end else begin
        tlbl2_6_flag_v <= _GEN_3486;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_v <= _GEN_1642;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_flag_v <= _GEN_1642;
    end else begin
      tlbl2_6_flag_v <= _GEN_2932;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_ppn <= _GEN_1658;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_ppn <= _GEN_1658;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_ppn <= _GEN_2733;
    end else begin
      tlbl2_6_ppn <= _GEN_1658;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_6_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_rmask <= _GEN_1674;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_rmask <= _GEN_1674;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_6_rmask <= _GEN_2749;
    end else begin
      tlbl2_6_rmask <= _GEN_1674;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_vpn <= _GEN_1499;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_vpn <= _GEN_1499;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_vpn <= _GEN_2574;
    end else begin
      tlbl2_7_vpn <= _GEN_1499;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_asid <= _GEN_1515;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_asid <= _GEN_1515;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_asid <= _GEN_2590;
    end else begin
      tlbl2_7_asid <= _GEN_1515;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_d <= _GEN_1531;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_d <= _GEN_1531;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_d <= _GEN_2606;
    end else begin
      tlbl2_7_flag_d <= _GEN_1531;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_g <= _GEN_1563;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_g <= _GEN_1563;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_g <= _GEN_2638;
    end else begin
      tlbl2_7_flag_g <= _GEN_1563;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_u <= _GEN_1579;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_u <= _GEN_1579;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_u <= _GEN_2654;
    end else begin
      tlbl2_7_flag_u <= _GEN_1579;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_x <= _GEN_1595;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_x <= _GEN_1595;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_x <= _GEN_2670;
    end else begin
      tlbl2_7_flag_x <= _GEN_1595;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_w <= _GEN_1611;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_w <= _GEN_1611;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_w <= _GEN_2686;
    end else begin
      tlbl2_7_flag_w <= _GEN_1611;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_r <= _GEN_1627;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_r <= _GEN_1627;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_r <= _GEN_2702;
    end else begin
      tlbl2_7_flag_r <= _GEN_1627;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_7_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_7_flag_v <= _GEN_3415;
      end else begin
        tlbl2_7_flag_v <= _GEN_3487;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_v <= _GEN_1643;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_flag_v <= _GEN_1643;
    end else begin
      tlbl2_7_flag_v <= _GEN_2933;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_ppn <= _GEN_1659;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_ppn <= _GEN_1659;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_ppn <= _GEN_2734;
    end else begin
      tlbl2_7_ppn <= _GEN_1659;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_7_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_rmask <= _GEN_1675;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_rmask <= _GEN_1675;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_7_rmask <= _GEN_2750;
    end else begin
      tlbl2_7_rmask <= _GEN_1675;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_vpn <= _GEN_1500;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_vpn <= _GEN_1500;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_vpn <= _GEN_2575;
    end else begin
      tlbl2_8_vpn <= _GEN_1500;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_asid <= _GEN_1516;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_asid <= _GEN_1516;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_asid <= _GEN_2591;
    end else begin
      tlbl2_8_asid <= _GEN_1516;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_d <= _GEN_1532;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_d <= _GEN_1532;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_d <= _GEN_2607;
    end else begin
      tlbl2_8_flag_d <= _GEN_1532;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_g <= _GEN_1564;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_g <= _GEN_1564;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_g <= _GEN_2639;
    end else begin
      tlbl2_8_flag_g <= _GEN_1564;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_u <= _GEN_1580;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_u <= _GEN_1580;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_u <= _GEN_2655;
    end else begin
      tlbl2_8_flag_u <= _GEN_1580;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_x <= _GEN_1596;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_x <= _GEN_1596;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_x <= _GEN_2671;
    end else begin
      tlbl2_8_flag_x <= _GEN_1596;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_w <= _GEN_1612;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_w <= _GEN_1612;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_w <= _GEN_2687;
    end else begin
      tlbl2_8_flag_w <= _GEN_1612;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_r <= _GEN_1628;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_r <= _GEN_1628;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_r <= _GEN_2703;
    end else begin
      tlbl2_8_flag_r <= _GEN_1628;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_8_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_8_flag_v <= _GEN_3416;
      end else begin
        tlbl2_8_flag_v <= _GEN_3488;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_v <= _GEN_1644;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_flag_v <= _GEN_1644;
    end else begin
      tlbl2_8_flag_v <= _GEN_2934;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_ppn <= _GEN_1660;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_ppn <= _GEN_1660;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_ppn <= _GEN_2735;
    end else begin
      tlbl2_8_ppn <= _GEN_1660;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_8_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_rmask <= _GEN_1676;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_rmask <= _GEN_1676;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_8_rmask <= _GEN_2751;
    end else begin
      tlbl2_8_rmask <= _GEN_1676;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_vpn <= _GEN_1501;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_vpn <= _GEN_1501;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_vpn <= _GEN_2576;
    end else begin
      tlbl2_9_vpn <= _GEN_1501;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_asid <= _GEN_1517;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_asid <= _GEN_1517;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_asid <= _GEN_2592;
    end else begin
      tlbl2_9_asid <= _GEN_1517;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_d <= _GEN_1533;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_d <= _GEN_1533;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_d <= _GEN_2608;
    end else begin
      tlbl2_9_flag_d <= _GEN_1533;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_g <= _GEN_1565;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_g <= _GEN_1565;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_g <= _GEN_2640;
    end else begin
      tlbl2_9_flag_g <= _GEN_1565;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_u <= _GEN_1581;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_u <= _GEN_1581;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_u <= _GEN_2656;
    end else begin
      tlbl2_9_flag_u <= _GEN_1581;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_x <= _GEN_1597;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_x <= _GEN_1597;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_x <= _GEN_2672;
    end else begin
      tlbl2_9_flag_x <= _GEN_1597;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_w <= _GEN_1613;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_w <= _GEN_1613;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_w <= _GEN_2688;
    end else begin
      tlbl2_9_flag_w <= _GEN_1613;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_r <= _GEN_1629;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_r <= _GEN_1629;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_r <= _GEN_2704;
    end else begin
      tlbl2_9_flag_r <= _GEN_1629;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_9_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_9_flag_v <= _GEN_3417;
      end else begin
        tlbl2_9_flag_v <= _GEN_3489;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_v <= _GEN_1645;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_flag_v <= _GEN_1645;
    end else begin
      tlbl2_9_flag_v <= _GEN_2935;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_ppn <= _GEN_1661;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_ppn <= _GEN_1661;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_ppn <= _GEN_2736;
    end else begin
      tlbl2_9_ppn <= _GEN_1661;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_9_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_rmask <= _GEN_1677;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_rmask <= _GEN_1677;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_9_rmask <= _GEN_2752;
    end else begin
      tlbl2_9_rmask <= _GEN_1677;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_vpn <= _GEN_1502;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_vpn <= _GEN_1502;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_vpn <= _GEN_2577;
    end else begin
      tlbl2_10_vpn <= _GEN_1502;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_asid <= _GEN_1518;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_asid <= _GEN_1518;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_asid <= _GEN_2593;
    end else begin
      tlbl2_10_asid <= _GEN_1518;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_d <= _GEN_1534;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_d <= _GEN_1534;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_d <= _GEN_2609;
    end else begin
      tlbl2_10_flag_d <= _GEN_1534;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_g <= _GEN_1566;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_g <= _GEN_1566;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_g <= _GEN_2641;
    end else begin
      tlbl2_10_flag_g <= _GEN_1566;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_u <= _GEN_1582;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_u <= _GEN_1582;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_u <= _GEN_2657;
    end else begin
      tlbl2_10_flag_u <= _GEN_1582;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_x <= _GEN_1598;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_x <= _GEN_1598;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_x <= _GEN_2673;
    end else begin
      tlbl2_10_flag_x <= _GEN_1598;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_w <= _GEN_1614;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_w <= _GEN_1614;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_w <= _GEN_2689;
    end else begin
      tlbl2_10_flag_w <= _GEN_1614;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_r <= _GEN_1630;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_r <= _GEN_1630;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_r <= _GEN_2705;
    end else begin
      tlbl2_10_flag_r <= _GEN_1630;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_10_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_10_flag_v <= _GEN_3418;
      end else begin
        tlbl2_10_flag_v <= _GEN_3490;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_v <= _GEN_1646;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_flag_v <= _GEN_1646;
    end else begin
      tlbl2_10_flag_v <= _GEN_2936;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_ppn <= _GEN_1662;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_ppn <= _GEN_1662;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_ppn <= _GEN_2737;
    end else begin
      tlbl2_10_ppn <= _GEN_1662;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_10_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_rmask <= _GEN_1678;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_rmask <= _GEN_1678;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_10_rmask <= _GEN_2753;
    end else begin
      tlbl2_10_rmask <= _GEN_1678;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_vpn <= _GEN_1503;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_vpn <= _GEN_1503;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_vpn <= _GEN_2578;
    end else begin
      tlbl2_11_vpn <= _GEN_1503;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_asid <= _GEN_1519;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_asid <= _GEN_1519;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_asid <= _GEN_2594;
    end else begin
      tlbl2_11_asid <= _GEN_1519;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_d <= _GEN_1535;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_d <= _GEN_1535;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_d <= _GEN_2610;
    end else begin
      tlbl2_11_flag_d <= _GEN_1535;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_g <= _GEN_1567;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_g <= _GEN_1567;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_g <= _GEN_2642;
    end else begin
      tlbl2_11_flag_g <= _GEN_1567;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_u <= _GEN_1583;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_u <= _GEN_1583;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_u <= _GEN_2658;
    end else begin
      tlbl2_11_flag_u <= _GEN_1583;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_x <= _GEN_1599;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_x <= _GEN_1599;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_x <= _GEN_2674;
    end else begin
      tlbl2_11_flag_x <= _GEN_1599;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_w <= _GEN_1615;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_w <= _GEN_1615;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_w <= _GEN_2690;
    end else begin
      tlbl2_11_flag_w <= _GEN_1615;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_r <= _GEN_1631;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_r <= _GEN_1631;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_r <= _GEN_2706;
    end else begin
      tlbl2_11_flag_r <= _GEN_1631;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_11_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_11_flag_v <= _GEN_3419;
      end else begin
        tlbl2_11_flag_v <= _GEN_3491;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_v <= _GEN_1647;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_flag_v <= _GEN_1647;
    end else begin
      tlbl2_11_flag_v <= _GEN_2937;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_ppn <= _GEN_1663;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_ppn <= _GEN_1663;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_ppn <= _GEN_2738;
    end else begin
      tlbl2_11_ppn <= _GEN_1663;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_11_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_rmask <= _GEN_1679;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_rmask <= _GEN_1679;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_11_rmask <= _GEN_2754;
    end else begin
      tlbl2_11_rmask <= _GEN_1679;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_vpn <= _GEN_1504;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_vpn <= _GEN_1504;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_vpn <= _GEN_2579;
    end else begin
      tlbl2_12_vpn <= _GEN_1504;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_asid <= _GEN_1520;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_asid <= _GEN_1520;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_asid <= _GEN_2595;
    end else begin
      tlbl2_12_asid <= _GEN_1520;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_d <= _GEN_1536;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_d <= _GEN_1536;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_d <= _GEN_2611;
    end else begin
      tlbl2_12_flag_d <= _GEN_1536;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_g <= _GEN_1568;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_g <= _GEN_1568;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_g <= _GEN_2643;
    end else begin
      tlbl2_12_flag_g <= _GEN_1568;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_u <= _GEN_1584;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_u <= _GEN_1584;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_u <= _GEN_2659;
    end else begin
      tlbl2_12_flag_u <= _GEN_1584;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_x <= _GEN_1600;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_x <= _GEN_1600;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_x <= _GEN_2675;
    end else begin
      tlbl2_12_flag_x <= _GEN_1600;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_w <= _GEN_1616;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_w <= _GEN_1616;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_w <= _GEN_2691;
    end else begin
      tlbl2_12_flag_w <= _GEN_1616;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_r <= _GEN_1632;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_r <= _GEN_1632;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_r <= _GEN_2707;
    end else begin
      tlbl2_12_flag_r <= _GEN_1632;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_12_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_12_flag_v <= _GEN_3420;
      end else begin
        tlbl2_12_flag_v <= _GEN_3492;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_v <= _GEN_1648;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_flag_v <= _GEN_1648;
    end else begin
      tlbl2_12_flag_v <= _GEN_2938;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_ppn <= _GEN_1664;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_ppn <= _GEN_1664;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_ppn <= _GEN_2739;
    end else begin
      tlbl2_12_ppn <= _GEN_1664;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_12_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_rmask <= _GEN_1680;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_rmask <= _GEN_1680;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_12_rmask <= _GEN_2755;
    end else begin
      tlbl2_12_rmask <= _GEN_1680;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_vpn <= _GEN_1505;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_vpn <= _GEN_1505;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_vpn <= _GEN_2580;
    end else begin
      tlbl2_13_vpn <= _GEN_1505;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_asid <= _GEN_1521;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_asid <= _GEN_1521;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_asid <= _GEN_2596;
    end else begin
      tlbl2_13_asid <= _GEN_1521;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_d <= _GEN_1537;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_d <= _GEN_1537;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_d <= _GEN_2612;
    end else begin
      tlbl2_13_flag_d <= _GEN_1537;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_g <= _GEN_1569;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_g <= _GEN_1569;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_g <= _GEN_2644;
    end else begin
      tlbl2_13_flag_g <= _GEN_1569;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_u <= _GEN_1585;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_u <= _GEN_1585;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_u <= _GEN_2660;
    end else begin
      tlbl2_13_flag_u <= _GEN_1585;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_x <= _GEN_1601;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_x <= _GEN_1601;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_x <= _GEN_2676;
    end else begin
      tlbl2_13_flag_x <= _GEN_1601;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_w <= _GEN_1617;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_w <= _GEN_1617;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_w <= _GEN_2692;
    end else begin
      tlbl2_13_flag_w <= _GEN_1617;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_r <= _GEN_1633;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_r <= _GEN_1633;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_r <= _GEN_2708;
    end else begin
      tlbl2_13_flag_r <= _GEN_1633;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_13_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_13_flag_v <= _GEN_3421;
      end else begin
        tlbl2_13_flag_v <= _GEN_3493;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_v <= _GEN_1649;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_flag_v <= _GEN_1649;
    end else begin
      tlbl2_13_flag_v <= _GEN_2939;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_ppn <= _GEN_1665;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_ppn <= _GEN_1665;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_ppn <= _GEN_2740;
    end else begin
      tlbl2_13_ppn <= _GEN_1665;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_13_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_rmask <= _GEN_1681;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_rmask <= _GEN_1681;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_13_rmask <= _GEN_2756;
    end else begin
      tlbl2_13_rmask <= _GEN_1681;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_vpn <= _GEN_1506;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_vpn <= _GEN_1506;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_vpn <= _GEN_2581;
    end else begin
      tlbl2_14_vpn <= _GEN_1506;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_asid <= _GEN_1522;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_asid <= _GEN_1522;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_asid <= _GEN_2597;
    end else begin
      tlbl2_14_asid <= _GEN_1522;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_d <= _GEN_1538;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_d <= _GEN_1538;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_d <= _GEN_2613;
    end else begin
      tlbl2_14_flag_d <= _GEN_1538;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_g <= _GEN_1570;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_g <= _GEN_1570;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_g <= _GEN_2645;
    end else begin
      tlbl2_14_flag_g <= _GEN_1570;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_u <= _GEN_1586;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_u <= _GEN_1586;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_u <= _GEN_2661;
    end else begin
      tlbl2_14_flag_u <= _GEN_1586;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_x <= _GEN_1602;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_x <= _GEN_1602;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_x <= _GEN_2677;
    end else begin
      tlbl2_14_flag_x <= _GEN_1602;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_w <= _GEN_1618;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_w <= _GEN_1618;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_w <= _GEN_2693;
    end else begin
      tlbl2_14_flag_w <= _GEN_1618;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_r <= _GEN_1634;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_r <= _GEN_1634;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_r <= _GEN_2709;
    end else begin
      tlbl2_14_flag_r <= _GEN_1634;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_14_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_14_flag_v <= _GEN_3422;
      end else begin
        tlbl2_14_flag_v <= _GEN_3494;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_v <= _GEN_1650;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_flag_v <= _GEN_1650;
    end else begin
      tlbl2_14_flag_v <= _GEN_2940;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_ppn <= _GEN_1666;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_ppn <= _GEN_1666;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_ppn <= _GEN_2741;
    end else begin
      tlbl2_14_ppn <= _GEN_1666;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_14_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_rmask <= _GEN_1682;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_rmask <= _GEN_1682;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_14_rmask <= _GEN_2757;
    end else begin
      tlbl2_14_rmask <= _GEN_1682;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_vpn <= 27'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_vpn <= _GEN_1507;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_vpn <= _GEN_1507;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_vpn <= _GEN_2582;
    end else begin
      tlbl2_15_vpn <= _GEN_1507;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_asid <= 16'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_asid <= _GEN_1523;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_asid <= _GEN_1523;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_asid <= _GEN_2598;
    end else begin
      tlbl2_15_asid <= _GEN_1523;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_d <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_d <= _GEN_1539;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_d <= _GEN_1539;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_d <= _GEN_2614;
    end else begin
      tlbl2_15_flag_d <= _GEN_1539;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_g <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_g <= _GEN_1571;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_g <= _GEN_1571;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_g <= _GEN_2646;
    end else begin
      tlbl2_15_flag_g <= _GEN_1571;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_u <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_u <= _GEN_1587;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_u <= _GEN_1587;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_u <= _GEN_2662;
    end else begin
      tlbl2_15_flag_u <= _GEN_1587;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_x <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_x <= _GEN_1603;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_x <= _GEN_1603;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_x <= _GEN_2678;
    end else begin
      tlbl2_15_flag_x <= _GEN_1603;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_w <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_w <= _GEN_1619;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_w <= _GEN_1619;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_w <= _GEN_2694;
    end else begin
      tlbl2_15_flag_w <= _GEN_1619;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_r <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_r <= _GEN_1635;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_r <= _GEN_1635;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_r <= _GEN_2710;
    end else begin
      tlbl2_15_flag_r <= _GEN_1635;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (io_sfence_vma_valid) begin // @[playground/src/cache/mmu/Tlb.scala 367:29]
      if (~(|src1) & ~(|src2)) begin // @[playground/src/cache/mmu/Tlb.scala 368:34]
        tlbl2_15_flag_v <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 373:25]
      end else if (_T_47 & _T_48) begin // @[playground/src/cache/mmu/Tlb.scala 375:39]
        tlbl2_15_flag_v <= _GEN_3423;
      end else begin
        tlbl2_15_flag_v <= _GEN_3495;
      end
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_v <= _GEN_1651;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_flag_v <= _GEN_1651;
    end else begin
      tlbl2_15_flag_v <= _GEN_2941;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_ppn <= 20'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_ppn <= _GEN_1667;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_ppn <= _GEN_1667;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_ppn <= _GEN_2742;
    end else begin
      tlbl2_15_ppn <= _GEN_1667;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 77:22]
      tlbl2_15_rmask <= 18'h0; // @[playground/src/cache/mmu/Tlb.scala 77:22]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_rmask <= _GEN_1683;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_rmask <= _GEN_1683;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      tlbl2_15_rmask <= _GEN_2758;
    end else begin
      tlbl2_15_rmask <= _GEN_1683;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 106:76]
      immu_state <= 2'h0; // @[playground/src/cache/mmu/Tlb.scala 106:76]
    end else if (2'h0 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (io_icache_en) begin // @[playground/src/cache/mmu/Tlb.scala 195:26]
        if (!(~ivm_enabled)) begin // @[playground/src/cache/mmu/Tlb.scala 199:28]
          immu_state <= _GEN_21;
        end
      end
    end else if (2'h1 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (|_T_9) begin // @[playground/src/cache/mmu/Tlb.scala 220:36]
        immu_state <= 2'h0; // @[playground/src/cache/mmu/Tlb.scala 221:20]
      end else begin
        immu_state <= _GEN_221;
      end
    end else if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      immu_state <= _GEN_844;
    end else begin
      immu_state <= _GEN_1056;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 107:76]
      dmmu_state <= 2'h0; // @[playground/src/cache/mmu/Tlb.scala 107:76]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (io_dcache_en) begin // @[playground/src/cache/mmu/Tlb.scala 268:26]
        if (!(~dvm_enabled)) begin // @[playground/src/cache/mmu/Tlb.scala 272:28]
          dmmu_state <= _GEN_1744;
        end
      end
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (|_T_40) begin // @[playground/src/cache/mmu/Tlb.scala 320:36]
        dmmu_state <= 2'h0; // @[playground/src/cache/mmu/Tlb.scala 321:20]
      end else begin
        dmmu_state <= _GEN_1944;
      end
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      dmmu_state <= _GEN_2565;
    end else begin
      dmmu_state <= _GEN_2777;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      replace_index_value <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      replace_index_value <= _GEN_1684;
    end else if (2'h1 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      replace_index_value <= _GEN_1684;
    end else if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      replace_index_value <= _GEN_2771;
    end else begin
      replace_index_value <= _GEN_1684;
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 112:30]
      ipage_fault <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 112:30]
    end else if (2'h0 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (io_icache_en) begin // @[playground/src/cache/mmu/Tlb.scala 195:26]
        if (~ivm_enabled) begin // @[playground/src/cache/mmu/Tlb.scala 199:28]
          ipage_fault <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 197:23]
        end else begin
          ipage_fault <= _GEN_20;
        end
      end
    end else if (!(2'h1 == immu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
      if (2'h2 == immu_state) begin // @[playground/src/cache/mmu/Tlb.scala 193:22]
        ipage_fault <= _GEN_845;
      end else begin
        ipage_fault <= _GEN_1054;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 113:30]
      dpage_fault <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 113:30]
    end else if (2'h0 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (io_dcache_en) begin // @[playground/src/cache/mmu/Tlb.scala 268:26]
        if (~dvm_enabled) begin // @[playground/src/cache/mmu/Tlb.scala 272:28]
          dpage_fault <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 270:23]
        end else begin
          dpage_fault <= _GEN_1743;
        end
      end
    end else if (!(2'h1 == dmmu_state)) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
      if (2'h2 == dmmu_state) begin // @[playground/src/cache/mmu/Tlb.scala 266:22]
        dpage_fault <= _GEN_2566;
      end else begin
        dpage_fault <= _GEN_2775;
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 120:28]
      ar_sel_lock <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 120:28]
    end else if (io_dcache_ptw_vpn_valid) begin // @[playground/src/cache/mmu/Tlb.scala 125:33]
      if (io_dcache_ptw_vpn_ready) begin // @[playground/src/cache/mmu/Tlb.scala 126:35]
        ar_sel_lock <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 127:19]
      end else begin
        ar_sel_lock <= 1'h1; // @[playground/src/cache/mmu/Tlb.scala 129:19]
      end
    end
    if (reset) begin // @[playground/src/cache/mmu/Tlb.scala 121:28]
      ar_sel_val <= 1'h0; // @[playground/src/cache/mmu/Tlb.scala 121:28]
    end else if (io_dcache_ptw_vpn_valid) begin // @[playground/src/cache/mmu/Tlb.scala 125:33]
      if (!(io_dcache_ptw_vpn_ready)) begin // @[playground/src/cache/mmu/Tlb.scala 126:35]
        if (!(ar_sel_lock)) begin // @[playground/src/cache/mmu/Tlb.scala 123:26]
          ar_sel_val <= req_ptw_0 & ~req_ptw_1;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  itlb_vpn = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  itlb_asid = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  itlb_flag_g = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  itlb_flag_u = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  itlb_flag_x = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  itlb_flag_v = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  itlb_ppn = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  itlb_rmask = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  dtlb_vpn = _RAND_8[26:0];
  _RAND_9 = {1{`RANDOM}};
  dtlb_asid = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  dtlb_flag_d = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dtlb_flag_g = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dtlb_flag_u = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  dtlb_flag_x = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dtlb_flag_w = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dtlb_flag_r = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dtlb_flag_v = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dtlb_ppn = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  dtlb_rmask = _RAND_18[17:0];
  _RAND_19 = {1{`RANDOM}};
  tlbl2_0_vpn = _RAND_19[26:0];
  _RAND_20 = {1{`RANDOM}};
  tlbl2_0_asid = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  tlbl2_0_flag_d = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  tlbl2_0_flag_g = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  tlbl2_0_flag_u = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  tlbl2_0_flag_x = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tlbl2_0_flag_w = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tlbl2_0_flag_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  tlbl2_0_flag_v = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  tlbl2_0_ppn = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  tlbl2_0_rmask = _RAND_29[17:0];
  _RAND_30 = {1{`RANDOM}};
  tlbl2_1_vpn = _RAND_30[26:0];
  _RAND_31 = {1{`RANDOM}};
  tlbl2_1_asid = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  tlbl2_1_flag_d = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlbl2_1_flag_g = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlbl2_1_flag_u = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tlbl2_1_flag_x = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tlbl2_1_flag_w = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  tlbl2_1_flag_r = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tlbl2_1_flag_v = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  tlbl2_1_ppn = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  tlbl2_1_rmask = _RAND_40[17:0];
  _RAND_41 = {1{`RANDOM}};
  tlbl2_2_vpn = _RAND_41[26:0];
  _RAND_42 = {1{`RANDOM}};
  tlbl2_2_asid = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  tlbl2_2_flag_d = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tlbl2_2_flag_g = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  tlbl2_2_flag_u = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  tlbl2_2_flag_x = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tlbl2_2_flag_w = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  tlbl2_2_flag_r = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  tlbl2_2_flag_v = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  tlbl2_2_ppn = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  tlbl2_2_rmask = _RAND_51[17:0];
  _RAND_52 = {1{`RANDOM}};
  tlbl2_3_vpn = _RAND_52[26:0];
  _RAND_53 = {1{`RANDOM}};
  tlbl2_3_asid = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  tlbl2_3_flag_d = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  tlbl2_3_flag_g = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  tlbl2_3_flag_u = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  tlbl2_3_flag_x = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  tlbl2_3_flag_w = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  tlbl2_3_flag_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  tlbl2_3_flag_v = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  tlbl2_3_ppn = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  tlbl2_3_rmask = _RAND_62[17:0];
  _RAND_63 = {1{`RANDOM}};
  tlbl2_4_vpn = _RAND_63[26:0];
  _RAND_64 = {1{`RANDOM}};
  tlbl2_4_asid = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  tlbl2_4_flag_d = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  tlbl2_4_flag_g = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  tlbl2_4_flag_u = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  tlbl2_4_flag_x = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  tlbl2_4_flag_w = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  tlbl2_4_flag_r = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tlbl2_4_flag_v = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  tlbl2_4_ppn = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  tlbl2_4_rmask = _RAND_73[17:0];
  _RAND_74 = {1{`RANDOM}};
  tlbl2_5_vpn = _RAND_74[26:0];
  _RAND_75 = {1{`RANDOM}};
  tlbl2_5_asid = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  tlbl2_5_flag_d = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  tlbl2_5_flag_g = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  tlbl2_5_flag_u = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  tlbl2_5_flag_x = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  tlbl2_5_flag_w = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  tlbl2_5_flag_r = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  tlbl2_5_flag_v = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  tlbl2_5_ppn = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  tlbl2_5_rmask = _RAND_84[17:0];
  _RAND_85 = {1{`RANDOM}};
  tlbl2_6_vpn = _RAND_85[26:0];
  _RAND_86 = {1{`RANDOM}};
  tlbl2_6_asid = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  tlbl2_6_flag_d = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  tlbl2_6_flag_g = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  tlbl2_6_flag_u = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  tlbl2_6_flag_x = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  tlbl2_6_flag_w = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  tlbl2_6_flag_r = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  tlbl2_6_flag_v = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  tlbl2_6_ppn = _RAND_94[19:0];
  _RAND_95 = {1{`RANDOM}};
  tlbl2_6_rmask = _RAND_95[17:0];
  _RAND_96 = {1{`RANDOM}};
  tlbl2_7_vpn = _RAND_96[26:0];
  _RAND_97 = {1{`RANDOM}};
  tlbl2_7_asid = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  tlbl2_7_flag_d = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  tlbl2_7_flag_g = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  tlbl2_7_flag_u = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  tlbl2_7_flag_x = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  tlbl2_7_flag_w = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  tlbl2_7_flag_r = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  tlbl2_7_flag_v = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  tlbl2_7_ppn = _RAND_105[19:0];
  _RAND_106 = {1{`RANDOM}};
  tlbl2_7_rmask = _RAND_106[17:0];
  _RAND_107 = {1{`RANDOM}};
  tlbl2_8_vpn = _RAND_107[26:0];
  _RAND_108 = {1{`RANDOM}};
  tlbl2_8_asid = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  tlbl2_8_flag_d = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  tlbl2_8_flag_g = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  tlbl2_8_flag_u = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  tlbl2_8_flag_x = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  tlbl2_8_flag_w = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  tlbl2_8_flag_r = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  tlbl2_8_flag_v = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  tlbl2_8_ppn = _RAND_116[19:0];
  _RAND_117 = {1{`RANDOM}};
  tlbl2_8_rmask = _RAND_117[17:0];
  _RAND_118 = {1{`RANDOM}};
  tlbl2_9_vpn = _RAND_118[26:0];
  _RAND_119 = {1{`RANDOM}};
  tlbl2_9_asid = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  tlbl2_9_flag_d = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  tlbl2_9_flag_g = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  tlbl2_9_flag_u = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  tlbl2_9_flag_x = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  tlbl2_9_flag_w = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  tlbl2_9_flag_r = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  tlbl2_9_flag_v = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  tlbl2_9_ppn = _RAND_127[19:0];
  _RAND_128 = {1{`RANDOM}};
  tlbl2_9_rmask = _RAND_128[17:0];
  _RAND_129 = {1{`RANDOM}};
  tlbl2_10_vpn = _RAND_129[26:0];
  _RAND_130 = {1{`RANDOM}};
  tlbl2_10_asid = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  tlbl2_10_flag_d = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  tlbl2_10_flag_g = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  tlbl2_10_flag_u = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  tlbl2_10_flag_x = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  tlbl2_10_flag_w = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  tlbl2_10_flag_r = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  tlbl2_10_flag_v = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  tlbl2_10_ppn = _RAND_138[19:0];
  _RAND_139 = {1{`RANDOM}};
  tlbl2_10_rmask = _RAND_139[17:0];
  _RAND_140 = {1{`RANDOM}};
  tlbl2_11_vpn = _RAND_140[26:0];
  _RAND_141 = {1{`RANDOM}};
  tlbl2_11_asid = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  tlbl2_11_flag_d = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  tlbl2_11_flag_g = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  tlbl2_11_flag_u = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  tlbl2_11_flag_x = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  tlbl2_11_flag_w = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  tlbl2_11_flag_r = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  tlbl2_11_flag_v = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  tlbl2_11_ppn = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  tlbl2_11_rmask = _RAND_150[17:0];
  _RAND_151 = {1{`RANDOM}};
  tlbl2_12_vpn = _RAND_151[26:0];
  _RAND_152 = {1{`RANDOM}};
  tlbl2_12_asid = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  tlbl2_12_flag_d = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  tlbl2_12_flag_g = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  tlbl2_12_flag_u = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tlbl2_12_flag_x = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tlbl2_12_flag_w = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  tlbl2_12_flag_r = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  tlbl2_12_flag_v = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  tlbl2_12_ppn = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  tlbl2_12_rmask = _RAND_161[17:0];
  _RAND_162 = {1{`RANDOM}};
  tlbl2_13_vpn = _RAND_162[26:0];
  _RAND_163 = {1{`RANDOM}};
  tlbl2_13_asid = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  tlbl2_13_flag_d = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  tlbl2_13_flag_g = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  tlbl2_13_flag_u = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  tlbl2_13_flag_x = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  tlbl2_13_flag_w = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  tlbl2_13_flag_r = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  tlbl2_13_flag_v = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  tlbl2_13_ppn = _RAND_171[19:0];
  _RAND_172 = {1{`RANDOM}};
  tlbl2_13_rmask = _RAND_172[17:0];
  _RAND_173 = {1{`RANDOM}};
  tlbl2_14_vpn = _RAND_173[26:0];
  _RAND_174 = {1{`RANDOM}};
  tlbl2_14_asid = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  tlbl2_14_flag_d = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  tlbl2_14_flag_g = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  tlbl2_14_flag_u = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  tlbl2_14_flag_x = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  tlbl2_14_flag_w = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  tlbl2_14_flag_r = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  tlbl2_14_flag_v = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  tlbl2_14_ppn = _RAND_182[19:0];
  _RAND_183 = {1{`RANDOM}};
  tlbl2_14_rmask = _RAND_183[17:0];
  _RAND_184 = {1{`RANDOM}};
  tlbl2_15_vpn = _RAND_184[26:0];
  _RAND_185 = {1{`RANDOM}};
  tlbl2_15_asid = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  tlbl2_15_flag_d = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  tlbl2_15_flag_g = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  tlbl2_15_flag_u = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  tlbl2_15_flag_x = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  tlbl2_15_flag_w = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  tlbl2_15_flag_r = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  tlbl2_15_flag_v = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  tlbl2_15_ppn = _RAND_193[19:0];
  _RAND_194 = {1{`RANDOM}};
  tlbl2_15_rmask = _RAND_194[17:0];
  _RAND_195 = {1{`RANDOM}};
  immu_state = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  dmmu_state = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  replace_index_value = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  ipage_fault = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dpage_fault = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ar_sel_lock = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ar_sel_val = _RAND_201[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_ext_int_ei, // @[playground/src/Core.scala 18:14]
  input         io_ext_int_ti, // @[playground/src/Core.scala 18:14]
  input         io_ext_int_si, // @[playground/src/Core.scala 18:14]
  output        io_inst_req, // @[playground/src/Core.scala 18:14]
  output        io_inst_complete_single_request, // @[playground/src/Core.scala 18:14]
  output [63:0] io_inst_addr_0, // @[playground/src/Core.scala 18:14]
  output [63:0] io_inst_addr_1, // @[playground/src/Core.scala 18:14]
  output        io_inst_fence_i, // @[playground/src/Core.scala 18:14]
  output        io_inst_dcache_stall, // @[playground/src/Core.scala 18:14]
  input  [63:0] io_inst_inst_0, // @[playground/src/Core.scala 18:14]
  input  [63:0] io_inst_inst_1, // @[playground/src/Core.scala 18:14]
  input         io_inst_inst_valid_0, // @[playground/src/Core.scala 18:14]
  input         io_inst_inst_valid_1, // @[playground/src/Core.scala 18:14]
  input         io_inst_access_fault, // @[playground/src/Core.scala 18:14]
  input         io_inst_page_fault, // @[playground/src/Core.scala 18:14]
  input         io_inst_addr_misaligned, // @[playground/src/Core.scala 18:14]
  input         io_inst_icache_stall, // @[playground/src/Core.scala 18:14]
  input         io_inst_tlb_en, // @[playground/src/Core.scala 18:14]
  input  [63:0] io_inst_tlb_vaddr, // @[playground/src/Core.scala 18:14]
  input         io_inst_tlb_complete_single_request, // @[playground/src/Core.scala 18:14]
  output        io_inst_tlb_uncached, // @[playground/src/Core.scala 18:14]
  output        io_inst_tlb_hit, // @[playground/src/Core.scala 18:14]
  output [19:0] io_inst_tlb_ptag, // @[playground/src/Core.scala 18:14]
  output [31:0] io_inst_tlb_paddr, // @[playground/src/Core.scala 18:14]
  output        io_inst_tlb_page_fault, // @[playground/src/Core.scala 18:14]
  output [63:0] io_data_exe_addr, // @[playground/src/Core.scala 18:14]
  output [63:0] io_data_addr, // @[playground/src/Core.scala 18:14]
  output [7:0]  io_data_rlen, // @[playground/src/Core.scala 18:14]
  output        io_data_en, // @[playground/src/Core.scala 18:14]
  output        io_data_wen, // @[playground/src/Core.scala 18:14]
  output [63:0] io_data_wdata, // @[playground/src/Core.scala 18:14]
  output        io_data_complete_single_request, // @[playground/src/Core.scala 18:14]
  output        io_data_fence_i, // @[playground/src/Core.scala 18:14]
  output [7:0]  io_data_wstrb, // @[playground/src/Core.scala 18:14]
  input  [63:0] io_data_rdata, // @[playground/src/Core.scala 18:14]
  input         io_data_access_fault, // @[playground/src/Core.scala 18:14]
  input         io_data_page_fault, // @[playground/src/Core.scala 18:14]
  input         io_data_dcache_ready, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_en, // @[playground/src/Core.scala 18:14]
  input  [63:0] io_data_tlb_vaddr, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_complete_single_request, // @[playground/src/Core.scala 18:14]
  output        io_data_tlb_uncached, // @[playground/src/Core.scala 18:14]
  output        io_data_tlb_hit, // @[playground/src/Core.scala 18:14]
  output [19:0] io_data_tlb_ptag, // @[playground/src/Core.scala 18:14]
  output [31:0] io_data_tlb_paddr, // @[playground/src/Core.scala 18:14]
  output        io_data_tlb_page_fault, // @[playground/src/Core.scala 18:14]
  input  [1:0]  io_data_tlb_access_type, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_vpn_ready, // @[playground/src/Core.scala 18:14]
  output        io_data_tlb_ptw_vpn_valid, // @[playground/src/Core.scala 18:14]
  output [26:0] io_data_tlb_ptw_vpn_bits, // @[playground/src/Core.scala 18:14]
  output [1:0]  io_data_tlb_ptw_access_type, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_valid, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_page_fault, // @[playground/src/Core.scala 18:14]
  input  [19:0] io_data_tlb_ptw_pte_bits_entry_ppn, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_d, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_g, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_u, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_x, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_w, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_r, // @[playground/src/Core.scala 18:14]
  input         io_data_tlb_ptw_pte_bits_entry_flag_v, // @[playground/src/Core.scala 18:14]
  input  [17:0] io_data_tlb_ptw_pte_bits_rmask, // @[playground/src/Core.scala 18:14]
  output [63:0] io_data_tlb_csr_satp, // @[playground/src/Core.scala 18:14]
  output [63:0] io_data_tlb_csr_mstatus, // @[playground/src/Core.scala 18:14]
  output [1:0]  io_data_tlb_csr_imode, // @[playground/src/Core.scala 18:14]
  output [1:0]  io_data_tlb_csr_dmode, // @[playground/src/Core.scala 18:14]
  output [63:0] io_debug_wb_pc, // @[playground/src/Core.scala 18:14]
  output        io_debug_wb_rf_wen, // @[playground/src/Core.scala 18:14]
  output [4:0]  io_debug_wb_rf_wnum, // @[playground/src/Core.scala 18:14]
  output [63:0] io_debug_wb_rf_wdata // @[playground/src/Core.scala 18:14]
);
  wire  Ctrl_io_cacheCtrl_iCache_stall; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_fetchUnit_allow_to_go; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_decodeUnit_inst0_src1_ren; // @[playground/src/Core.scala 25:30]
  wire [4:0] Ctrl_io_decodeUnit_inst0_src1_raddr; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_decodeUnit_inst0_src2_ren; // @[playground/src/Core.scala 25:30]
  wire [4:0] Ctrl_io_decodeUnit_inst0_src2_raddr; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_decodeUnit_branch; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_decodeUnit_allow_to_go; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_decodeUnit_do_flush; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_inst_0_is_load; // @[playground/src/Core.scala 25:30]
  wire [4:0] Ctrl_io_executeUnit_inst_0_reg_waddr; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_inst_1_is_load; // @[playground/src/Core.scala 25:30]
  wire [4:0] Ctrl_io_executeUnit_inst_1_reg_waddr; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_flush; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_allow_to_go; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_do_flush; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_fu_allow_to_go; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_executeUnit_fu_stall; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_memoryUnit_flush; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_memoryUnit_mem_stall; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_memoryUnit_allow_to_go; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_memoryUnit_do_flush; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_memoryUnit_complete_single_request; // @[playground/src/Core.scala 25:30]
  wire  Ctrl_io_writeBackUnit_allow_to_go; // @[playground/src/Core.scala 25:30]
  wire  FetchUnit_clock; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_reset; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_io_memory_flush; // @[playground/src/Core.scala 26:30]
  wire [63:0] FetchUnit_io_memory_target; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_io_decode_branch; // @[playground/src/Core.scala 26:30]
  wire [63:0] FetchUnit_io_decode_target; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_io_execute_flush; // @[playground/src/Core.scala 26:30]
  wire [63:0] FetchUnit_io_execute_target; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_io_instFifo_full; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_io_iCache_inst_valid_0; // @[playground/src/Core.scala 26:30]
  wire  FetchUnit_io_iCache_inst_valid_1; // @[playground/src/Core.scala 26:30]
  wire [63:0] FetchUnit_io_iCache_pc; // @[playground/src/Core.scala 26:30]
  wire [63:0] FetchUnit_io_iCache_pc_next; // @[playground/src/Core.scala 26:30]
  wire  BranchPredictorUnit_clock; // @[playground/src/Core.scala 27:30]
  wire  BranchPredictorUnit_reset; // @[playground/src/Core.scala 27:30]
  wire [63:0] BranchPredictorUnit_io_decode_pc; // @[playground/src/Core.scala 27:30]
  wire  BranchPredictorUnit_io_decode_info_valid; // @[playground/src/Core.scala 27:30]
  wire [2:0] BranchPredictorUnit_io_decode_info_fusel; // @[playground/src/Core.scala 27:30]
  wire [6:0] BranchPredictorUnit_io_decode_info_op; // @[playground/src/Core.scala 27:30]
  wire [63:0] BranchPredictorUnit_io_decode_info_imm; // @[playground/src/Core.scala 27:30]
  wire [5:0] BranchPredictorUnit_io_decode_pht_index; // @[playground/src/Core.scala 27:30]
  wire  BranchPredictorUnit_io_decode_branch_inst; // @[playground/src/Core.scala 27:30]
  wire  BranchPredictorUnit_io_decode_branch; // @[playground/src/Core.scala 27:30]
  wire [63:0] BranchPredictorUnit_io_decode_target; // @[playground/src/Core.scala 27:30]
  wire [5:0] BranchPredictorUnit_io_decode_update_pht_index; // @[playground/src/Core.scala 27:30]
  wire [63:0] BranchPredictorUnit_io_instBuffer_pc_0; // @[playground/src/Core.scala 27:30]
  wire [63:0] BranchPredictorUnit_io_instBuffer_pc_1; // @[playground/src/Core.scala 27:30]
  wire [5:0] BranchPredictorUnit_io_instBuffer_pht_index_0; // @[playground/src/Core.scala 27:30]
  wire [5:0] BranchPredictorUnit_io_instBuffer_pht_index_1; // @[playground/src/Core.scala 27:30]
  wire [63:0] BranchPredictorUnit_io_execute_pc; // @[playground/src/Core.scala 27:30]
  wire [5:0] BranchPredictorUnit_io_execute_update_pht_index; // @[playground/src/Core.scala 27:30]
  wire  BranchPredictorUnit_io_execute_branch_inst; // @[playground/src/Core.scala 27:30]
  wire  BranchPredictorUnit_io_execute_branch; // @[playground/src/Core.scala 27:30]
  wire  InstFifo_clock; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_reset; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_do_flush; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_wen_0; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_wen_1; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_write_0_inst; // @[playground/src/Core.scala 28:30]
  wire [5:0] InstFifo_io_write_0_pht_index; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_write_0_addr_misaligned; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_write_0_access_fault; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_write_0_page_fault; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_write_0_pc; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_write_1_inst; // @[playground/src/Core.scala 28:30]
  wire [5:0] InstFifo_io_write_1_pht_index; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_write_1_addr_misaligned; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_write_1_access_fault; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_write_1_page_fault; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_write_1_pc; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_full; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_allow_to_go_0; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_allow_to_go_1; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_decoderUint_inst_0_inst; // @[playground/src/Core.scala 28:30]
  wire [5:0] InstFifo_io_decoderUint_inst_0_pht_index; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_inst_0_addr_misaligned; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_inst_0_access_fault; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_inst_0_page_fault; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_decoderUint_inst_0_pc; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_decoderUint_inst_1_inst; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_inst_1_addr_misaligned; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_inst_1_access_fault; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_inst_1_page_fault; // @[playground/src/Core.scala 28:30]
  wire [63:0] InstFifo_io_decoderUint_inst_1_pc; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_info_empty; // @[playground/src/Core.scala 28:30]
  wire  InstFifo_io_decoderUint_info_almost_empty; // @[playground/src/Core.scala 28:30]
  wire  DecodeUnit_io_instFifo_allow_to_go_0; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_allow_to_go_1; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_instFifo_inst_0_inst; // @[playground/src/Core.scala 29:30]
  wire [5:0] DecodeUnit_io_instFifo_inst_0_pht_index; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_inst_0_addr_misaligned; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_inst_0_access_fault; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_inst_0_page_fault; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_instFifo_inst_0_pc; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_instFifo_inst_1_inst; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_inst_1_addr_misaligned; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_inst_1_access_fault; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_inst_1_page_fault; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_instFifo_inst_1_pc; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_info_empty; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_instFifo_info_almost_empty; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_regfile_0_src1_raddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_regfile_0_src1_rdata; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_regfile_0_src2_raddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_regfile_0_src2_rdata; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_regfile_1_src1_raddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_regfile_1_src1_rdata; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_regfile_1_src2_raddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_regfile_1_src2_rdata; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_forward_0_exe_wen; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_forward_0_exe_waddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_forward_0_exe_wdata; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_forward_0_is_load; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_forward_0_mem_wen; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_forward_0_mem_waddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_forward_0_mem_wdata; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_forward_1_exe_wen; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_forward_1_exe_waddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_forward_1_exe_wdata; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_forward_1_is_load; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_forward_1_mem_wen; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_forward_1_mem_waddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_forward_1_mem_wdata; // @[playground/src/Core.scala 29:30]
  wire [1:0] DecodeUnit_io_csr_mode; // @[playground/src/Core.scala 29:30]
  wire [11:0] DecodeUnit_io_csr_interrupt; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_fetchUnit_branch; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_fetchUnit_target; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_bpu_pc; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_bpu_info_valid; // @[playground/src/Core.scala 29:30]
  wire [2:0] DecodeUnit_io_bpu_info_fusel; // @[playground/src/Core.scala 29:30]
  wire [6:0] DecodeUnit_io_bpu_info_op; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_bpu_info_imm; // @[playground/src/Core.scala 29:30]
  wire [5:0] DecodeUnit_io_bpu_pht_index; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_bpu_branch_inst; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_bpu_branch; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_bpu_target; // @[playground/src/Core.scala 29:30]
  wire [5:0] DecodeUnit_io_bpu_update_pht_index; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_pc; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_info_valid; // @[playground/src/Core.scala 29:30]
  wire [2:0] DecodeUnit_io_executeStage_inst_0_info_fusel; // @[playground/src/Core.scala 29:30]
  wire [6:0] DecodeUnit_io_executeStage_inst_0_info_op; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_executeStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_info_imm; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_info_inst; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_src_info_src1_data; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_src_info_src2_data; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_pc; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_info_valid; // @[playground/src/Core.scala 29:30]
  wire [2:0] DecodeUnit_io_executeStage_inst_1_info_fusel; // @[playground/src/Core.scala 29:30]
  wire [6:0] DecodeUnit_io_executeStage_inst_1_info_op; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_executeStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_info_imm; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_info_inst; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_src_info_src1_data; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_src_info_src2_data; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_jump_branch_info_jump_regiser; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_jump_branch_info_branch_inst; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_executeStage_jump_branch_info_pred_branch; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_jump_branch_info_branch_target; // @[playground/src/Core.scala 29:30]
  wire [63:0] DecodeUnit_io_executeStage_jump_branch_info_update_pht_index; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_ctrl_inst0_src1_ren; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_ctrl_inst0_src1_raddr; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_ctrl_inst0_src2_ren; // @[playground/src/Core.scala 29:30]
  wire [4:0] DecodeUnit_io_ctrl_inst0_src2_raddr; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_ctrl_branch; // @[playground/src/Core.scala 29:30]
  wire  DecodeUnit_io_ctrl_allow_to_go; // @[playground/src/Core.scala 29:30]
  wire  ARegFile_clock; // @[playground/src/Core.scala 30:30]
  wire  ARegFile_reset; // @[playground/src/Core.scala 30:30]
  wire [4:0] ARegFile_io_read_0_src1_raddr; // @[playground/src/Core.scala 30:30]
  wire [63:0] ARegFile_io_read_0_src1_rdata; // @[playground/src/Core.scala 30:30]
  wire [4:0] ARegFile_io_read_0_src2_raddr; // @[playground/src/Core.scala 30:30]
  wire [63:0] ARegFile_io_read_0_src2_rdata; // @[playground/src/Core.scala 30:30]
  wire [4:0] ARegFile_io_read_1_src1_raddr; // @[playground/src/Core.scala 30:30]
  wire [63:0] ARegFile_io_read_1_src1_rdata; // @[playground/src/Core.scala 30:30]
  wire [4:0] ARegFile_io_read_1_src2_raddr; // @[playground/src/Core.scala 30:30]
  wire [63:0] ARegFile_io_read_1_src2_rdata; // @[playground/src/Core.scala 30:30]
  wire  ARegFile_io_write_0_wen; // @[playground/src/Core.scala 30:30]
  wire [4:0] ARegFile_io_write_0_waddr; // @[playground/src/Core.scala 30:30]
  wire [63:0] ARegFile_io_write_0_wdata; // @[playground/src/Core.scala 30:30]
  wire  ARegFile_io_write_1_wen; // @[playground/src/Core.scala 30:30]
  wire [4:0] ARegFile_io_write_1_waddr; // @[playground/src/Core.scala 30:30]
  wire [63:0] ARegFile_io_write_1_wdata; // @[playground/src/Core.scala 30:30]
  wire  ExecuteStage_clock; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_reset; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_ctrl_allow_to_go_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_ctrl_allow_to_go_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_ctrl_clear_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_ctrl_clear_1; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_pc; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_info_valid; // @[playground/src/Core.scala 31:30]
  wire [2:0] ExecuteStage_io_decodeUnit_inst_0_info_fusel; // @[playground/src/Core.scala 31:30]
  wire [6:0] ExecuteStage_io_decodeUnit_inst_0_info_op; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 31:30]
  wire [4:0] ExecuteStage_io_decodeUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_info_imm; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_info_inst; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_src_info_src1_data; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_src_info_src2_data; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_ex_tval_0; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_ex_tval_1; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_ex_tval_2; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_0_ex_tval_12; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_pc; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_info_valid; // @[playground/src/Core.scala 31:30]
  wire [2:0] ExecuteStage_io_decodeUnit_inst_1_info_fusel; // @[playground/src/Core.scala 31:30]
  wire [6:0] ExecuteStage_io_decodeUnit_inst_1_info_op; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 31:30]
  wire [4:0] ExecuteStage_io_decodeUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_info_imm; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_info_inst; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_src_info_src1_data; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_src_info_src2_data; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_ex_tval_0; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_ex_tval_1; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_ex_tval_2; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_inst_1_ex_tval_12; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_jump_branch_info_jump_regiser; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_jump_branch_info_branch_inst; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_decodeUnit_jump_branch_info_pred_branch; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_jump_branch_info_branch_target; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_decodeUnit_jump_branch_info_update_pht_index; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_pc; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_info_valid; // @[playground/src/Core.scala 31:30]
  wire [2:0] ExecuteStage_io_executeUnit_inst_0_info_fusel; // @[playground/src/Core.scala 31:30]
  wire [6:0] ExecuteStage_io_executeUnit_inst_0_info_op; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 31:30]
  wire [4:0] ExecuteStage_io_executeUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_info_imm; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_info_inst; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_src_info_src1_data; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_src_info_src2_data; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_ex_tval_0; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_ex_tval_1; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_ex_tval_2; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_0_ex_tval_12; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_pc; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_info_valid; // @[playground/src/Core.scala 31:30]
  wire [2:0] ExecuteStage_io_executeUnit_inst_1_info_fusel; // @[playground/src/Core.scala 31:30]
  wire [6:0] ExecuteStage_io_executeUnit_inst_1_info_op; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 31:30]
  wire [4:0] ExecuteStage_io_executeUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_info_imm; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_info_inst; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_src_info_src1_data; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_src_info_src2_data; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_ex_tval_0; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_ex_tval_1; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_ex_tval_2; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_inst_1_ex_tval_12; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_jump_branch_info_jump_regiser; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_jump_branch_info_branch_inst; // @[playground/src/Core.scala 31:30]
  wire  ExecuteStage_io_executeUnit_jump_branch_info_pred_branch; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_jump_branch_info_branch_target; // @[playground/src/Core.scala 31:30]
  wire [63:0] ExecuteStage_io_executeUnit_jump_branch_info_update_pht_index; // @[playground/src/Core.scala 31:30]
  wire  ExecuteUnit_clock; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_reset; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_ctrl_inst_0_is_load; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_ctrl_inst_0_reg_waddr; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_ctrl_inst_1_is_load; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_ctrl_inst_1_reg_waddr; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_ctrl_flush; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_ctrl_allow_to_go; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_ctrl_fu_allow_to_go; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_ctrl_fu_stall; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_pc; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_info_valid; // @[playground/src/Core.scala 32:30]
  wire [2:0] ExecuteUnit_io_executeStage_inst_0_info_fusel; // @[playground/src/Core.scala 32:30]
  wire [6:0] ExecuteUnit_io_executeStage_inst_0_info_op; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_executeStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_info_imm; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_info_inst; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_src_info_src1_data; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_src_info_src2_data; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_pc; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_info_valid; // @[playground/src/Core.scala 32:30]
  wire [2:0] ExecuteUnit_io_executeStage_inst_1_info_fusel; // @[playground/src/Core.scala 32:30]
  wire [6:0] ExecuteUnit_io_executeStage_inst_1_info_op; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_executeStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_info_imm; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_info_inst; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_src_info_src1_data; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_src_info_src2_data; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_jump_branch_info_jump_regiser; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_jump_branch_info_branch_inst; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_executeStage_jump_branch_info_pred_branch; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_jump_branch_info_branch_target; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_executeStage_jump_branch_info_update_pht_index; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_valid; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_in_pc; // @[playground/src/Core.scala 32:30]
  wire [6:0] ExecuteUnit_io_csr_in_info_op; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_in_info_inst; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_in_src_info_src1_data; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_11; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_exception_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_4; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_5; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_6; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_7; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_10; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_in_ex_interrupt_11; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_in_ex_tval_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_in_ex_tval_12; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_out_rdata; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_11; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_exception_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_4; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_5; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_6; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_7; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_10; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_ex_interrupt_11; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_out_ex_tval_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_out_ex_tval_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_out_ex_tval_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_csr_out_flush; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_csr_out_target; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_bpu_pc; // @[playground/src/Core.scala 32:30]
  wire [5:0] ExecuteUnit_io_bpu_update_pht_index; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_bpu_branch_inst; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_bpu_branch; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_fetchUnit_flush; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_fetchUnit_target; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_decodeUnit_forward_0_exe_wen; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_decodeUnit_forward_0_exe_waddr; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_decodeUnit_forward_0_exe_wdata; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_decodeUnit_forward_0_is_load; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_decodeUnit_forward_1_exe_wen; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_decodeUnit_forward_1_exe_waddr; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_decodeUnit_forward_1_exe_wdata; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_decodeUnit_forward_1_is_load; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_pc; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_info_valid; // @[playground/src/Core.scala 32:30]
  wire [2:0] ExecuteUnit_io_memoryStage_inst_0_info_fusel; // @[playground/src/Core.scala 32:30]
  wire [6:0] ExecuteUnit_io_memoryStage_inst_0_info_op; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_memoryStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_info_imm; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_info_inst; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_4; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_src_info_src1_data; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_src_info_src2_data; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_pc; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_info_valid; // @[playground/src/Core.scala 32:30]
  wire [2:0] ExecuteUnit_io_memoryStage_inst_1_info_fusel; // @[playground/src/Core.scala 32:30]
  wire [6:0] ExecuteUnit_io_memoryStage_inst_1_info_op; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 32:30]
  wire [4:0] ExecuteUnit_io_memoryStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_info_imm; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_info_inst; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_4; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_src_info_src1_data; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_src_info_src2_data; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 32:30]
  wire  ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_memoryStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 32:30]
  wire [63:0] ExecuteUnit_io_dataMemory_addr; // @[playground/src/Core.scala 32:30]
  wire  Csr_clock; // @[playground/src/Core.scala 33:30]
  wire  Csr_reset; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_ext_int_ei; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_ext_int_ti; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_ext_int_si; // @[playground/src/Core.scala 33:30]
  wire [1:0] Csr_io_decodeUnit_mode; // @[playground/src/Core.scala 33:30]
  wire [11:0] Csr_io_decodeUnit_interrupt; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_valid; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_in_pc; // @[playground/src/Core.scala 33:30]
  wire [6:0] Csr_io_executeUnit_in_info_op; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_in_info_inst; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_in_src_info_src1_data; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_1; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_2; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_3; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_8; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_9; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_11; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_exception_12; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_0; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_1; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_2; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_3; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_4; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_5; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_6; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_7; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_8; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_9; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_10; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_in_ex_interrupt_11; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_in_ex_tval_1; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_in_ex_tval_12; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_out_rdata; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_1; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_2; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_3; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_8; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_9; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_11; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_exception_12; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_0; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_1; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_2; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_3; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_4; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_5; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_6; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_7; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_8; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_9; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_10; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_ex_interrupt_11; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_out_ex_tval_1; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_out_ex_tval_2; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_out_ex_tval_12; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_executeUnit_out_flush; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_executeUnit_out_target; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_pc; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_0; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_1; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_2; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_3; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_4; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_5; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_6; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_7; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_8; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_9; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_10; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_11; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_12; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_13; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_14; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_exception_15; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_0; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_1; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_2; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_3; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_4; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_5; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_6; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_7; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_8; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_9; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_10; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_ex_interrupt_11; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_0; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_1; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_2; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_3; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_4; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_5; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_6; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_7; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_8; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_9; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_10; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_11; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_12; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_13; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_14; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_ex_tval_15; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_info_valid; // @[playground/src/Core.scala 33:30]
  wire [2:0] Csr_io_memoryUnit_in_info_fusel; // @[playground/src/Core.scala 33:30]
  wire [6:0] Csr_io_memoryUnit_in_info_op; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_lr_wen; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_in_lr_wbit; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_in_lr_waddr; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_out_flush; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_out_target; // @[playground/src/Core.scala 33:30]
  wire  Csr_io_memoryUnit_out_lr; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_memoryUnit_out_lr_addr; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_tlb_satp; // @[playground/src/Core.scala 33:30]
  wire [63:0] Csr_io_tlb_mstatus; // @[playground/src/Core.scala 33:30]
  wire [1:0] Csr_io_tlb_imode; // @[playground/src/Core.scala 33:30]
  wire [1:0] Csr_io_tlb_dmode; // @[playground/src/Core.scala 33:30]
  wire  MemoryStage_clock; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_reset; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_ctrl_allow_to_go; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_ctrl_clear; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_pc; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_info_valid; // @[playground/src/Core.scala 34:30]
  wire [2:0] MemoryStage_io_executeUnit_inst_0_info_fusel; // @[playground/src/Core.scala 34:30]
  wire [6:0] MemoryStage_io_executeUnit_inst_0_info_op; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 34:30]
  wire [4:0] MemoryStage_io_executeUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_info_imm; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_info_inst; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_src_info_src1_data; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_src_info_src2_data; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_ex_tval_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_ex_tval_1; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_ex_tval_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_0_ex_tval_12; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_pc; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_info_valid; // @[playground/src/Core.scala 34:30]
  wire [2:0] MemoryStage_io_executeUnit_inst_1_info_fusel; // @[playground/src/Core.scala 34:30]
  wire [6:0] MemoryStage_io_executeUnit_inst_1_info_op; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 34:30]
  wire [4:0] MemoryStage_io_executeUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_info_imm; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_info_inst; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_src_info_src1_data; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_src_info_src2_data; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_executeUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_ex_tval_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_ex_tval_1; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_ex_tval_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_executeUnit_inst_1_ex_tval_12; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_pc; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_info_valid; // @[playground/src/Core.scala 34:30]
  wire [2:0] MemoryStage_io_memoryUnit_inst_0_info_fusel; // @[playground/src/Core.scala 34:30]
  wire [6:0] MemoryStage_io_memoryUnit_inst_0_info_op; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 34:30]
  wire [4:0] MemoryStage_io_memoryUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_info_imm; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_info_inst; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_src_info_src1_data; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_src_info_src2_data; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_ex_tval_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_ex_tval_1; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_ex_tval_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_0_ex_tval_12; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_pc; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_info_valid; // @[playground/src/Core.scala 34:30]
  wire [2:0] MemoryStage_io_memoryUnit_inst_1_info_fusel; // @[playground/src/Core.scala 34:30]
  wire [6:0] MemoryStage_io_memoryUnit_inst_1_info_op; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 34:30]
  wire [4:0] MemoryStage_io_memoryUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_info_imm; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_info_inst; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_src_info_src1_data; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_src_info_src2_data; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 34:30]
  wire  MemoryStage_io_memoryUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_ex_tval_0; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_ex_tval_1; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_ex_tval_2; // @[playground/src/Core.scala 34:30]
  wire [63:0] MemoryStage_io_memoryUnit_inst_1_ex_tval_12; // @[playground/src/Core.scala 34:30]
  wire  MemoryUnit_clock; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_reset; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_ctrl_flush; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_ctrl_mem_stall; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_ctrl_allow_to_go; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_ctrl_fence_i; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_ctrl_complete_single_request; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_ctrl_sfence_vma_valid; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_ctrl_sfence_vma_src_info_src1_data; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_ctrl_sfence_vma_src_info_src2_data; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_pc; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_info_valid; // @[playground/src/Core.scala 35:30]
  wire [2:0] MemoryUnit_io_memoryStage_inst_0_info_fusel; // @[playground/src/Core.scala 35:30]
  wire [6:0] MemoryUnit_io_memoryStage_inst_0_info_op; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 35:30]
  wire [4:0] MemoryUnit_io_memoryStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_info_imm; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_info_inst; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_src_info_src1_data; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_src_info_src2_data; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_pc; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_info_valid; // @[playground/src/Core.scala 35:30]
  wire [2:0] MemoryUnit_io_memoryStage_inst_1_info_fusel; // @[playground/src/Core.scala 35:30]
  wire [6:0] MemoryUnit_io_memoryStage_inst_1_info_op; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 35:30]
  wire [4:0] MemoryUnit_io_memoryStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_info_imm; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_info_inst; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_src_info_src1_data; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_src_info_src2_data; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_memoryStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_memoryStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_fetchUnit_flush; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_fetchUnit_target; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_decodeUnit_0_wen; // @[playground/src/Core.scala 35:30]
  wire [4:0] MemoryUnit_io_decodeUnit_0_waddr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_decodeUnit_0_wdata; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_decodeUnit_1_wen; // @[playground/src/Core.scala 35:30]
  wire [4:0] MemoryUnit_io_decodeUnit_1_waddr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_decodeUnit_1_wdata; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_pc; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_11; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_12; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_13; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_14; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_exception_15; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_ex_interrupt_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_4; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_5; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_6; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_7; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_8; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_9; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_10; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_12; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_13; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_14; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_ex_tval_15; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_info_valid; // @[playground/src/Core.scala 35:30]
  wire [2:0] MemoryUnit_io_csr_in_info_fusel; // @[playground/src/Core.scala 35:30]
  wire [6:0] MemoryUnit_io_csr_in_info_op; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_lr_wen; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_in_lr_wbit; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_in_lr_waddr; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_out_flush; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_out_target; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_csr_out_lr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_csr_out_lr_addr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_pc; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_info_valid; // @[playground/src/Core.scala 35:30]
  wire [2:0] MemoryUnit_io_writeBackStage_inst_0_info_fusel; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 35:30]
  wire [4:0] MemoryUnit_io_writeBackStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_4; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_13; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_14; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_exception_15; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_4; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_5; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_6; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_7; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_8; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_9; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_10; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_13; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_14; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_0_ex_tval_15; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_pc; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_info_valid; // @[playground/src/Core.scala 35:30]
  wire [2:0] MemoryUnit_io_writeBackStage_inst_1_info_fusel; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 35:30]
  wire [4:0] MemoryUnit_io_writeBackStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_4; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_13; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_14; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_exception_15; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_3; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_4; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_5; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_6; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_7; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_8; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_9; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_10; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_11; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_13; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_14; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_writeBackStage_inst_1_ex_tval_15; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_dataMemory_in_access_fault; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_dataMemory_in_page_fault; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_dataMemory_in_ready; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_dataMemory_in_rdata; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_dataMemory_out_en; // @[playground/src/Core.scala 35:30]
  wire [7:0] MemoryUnit_io_dataMemory_out_rlen; // @[playground/src/Core.scala 35:30]
  wire  MemoryUnit_io_dataMemory_out_wen; // @[playground/src/Core.scala 35:30]
  wire [7:0] MemoryUnit_io_dataMemory_out_wstrb; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_dataMemory_out_addr; // @[playground/src/Core.scala 35:30]
  wire [63:0] MemoryUnit_io_dataMemory_out_wdata; // @[playground/src/Core.scala 35:30]
  wire  WriteBackStage_clock; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_reset; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_ctrl_allow_to_go; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_0_pc; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_info_valid; // @[playground/src/Core.scala 36:30]
  wire [2:0] WriteBackStage_io_memoryUnit_inst_0_info_fusel; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 36:30]
  wire [4:0] WriteBackStage_io_memoryUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_1; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_13; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_exception_15; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_1_pc; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_info_valid; // @[playground/src/Core.scala 36:30]
  wire [2:0] WriteBackStage_io_memoryUnit_inst_1_info_fusel; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 36:30]
  wire [4:0] WriteBackStage_io_memoryUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_1; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_13; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_exception_15; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_0_pc; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_info_valid; // @[playground/src/Core.scala 36:30]
  wire [2:0] WriteBackStage_io_writeBackUnit_inst_0_info_fusel; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 36:30]
  wire [4:0] WriteBackStage_io_writeBackUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_1; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_13; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_exception_15; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_1_pc; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_info_valid; // @[playground/src/Core.scala 36:30]
  wire [2:0] WriteBackStage_io_writeBackUnit_inst_1_info_fusel; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 36:30]
  wire [4:0] WriteBackStage_io_writeBackUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_1; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 36:30]
  wire [63:0] WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_13; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_exception_15; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 36:30]
  wire  WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 36:30]
  wire  WriteBackUnit_clock; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_ctrl_allow_to_go; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_0_pc; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_info_valid; // @[playground/src/Core.scala 37:30]
  wire [2:0] WriteBackUnit_io_writeBackStage_inst_0_info_fusel; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 37:30]
  wire [4:0] WriteBackUnit_io_writeBackStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_1; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_4; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_5; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_6; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_7; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_13; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_exception_15; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_1_pc; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_info_valid; // @[playground/src/Core.scala 37:30]
  wire [2:0] WriteBackUnit_io_writeBackStage_inst_1_info_fusel; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 37:30]
  wire [4:0] WriteBackUnit_io_writeBackStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_1; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_4; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_5; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_6; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_7; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_13; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_exception_15; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_regfile_0_wen; // @[playground/src/Core.scala 37:30]
  wire [4:0] WriteBackUnit_io_regfile_0_waddr; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_regfile_0_wdata; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_regfile_1_wen; // @[playground/src/Core.scala 37:30]
  wire [4:0] WriteBackUnit_io_regfile_1_waddr; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_regfile_1_wdata; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_debug_wb_pc; // @[playground/src/Core.scala 37:30]
  wire  WriteBackUnit_io_debug_wb_rf_wen; // @[playground/src/Core.scala 37:30]
  wire [4:0] WriteBackUnit_io_debug_wb_rf_wnum; // @[playground/src/Core.scala 37:30]
  wire [63:0] WriteBackUnit_io_debug_wb_rf_wdata; // @[playground/src/Core.scala 37:30]
  wire  Tlb_clock; // @[playground/src/Core.scala 38:30]
  wire  Tlb_reset; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_icache_en; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_icache_vaddr; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_icache_complete_single_request; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_icache_uncached; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_icache_hit; // @[playground/src/Core.scala 38:30]
  wire [19:0] Tlb_io_icache_ptag; // @[playground/src/Core.scala 38:30]
  wire [31:0] Tlb_io_icache_paddr; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_icache_page_fault; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_en; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_dcache_vaddr; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_complete_single_request; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_uncached; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_hit; // @[playground/src/Core.scala 38:30]
  wire [19:0] Tlb_io_dcache_ptag; // @[playground/src/Core.scala 38:30]
  wire [31:0] Tlb_io_dcache_paddr; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_page_fault; // @[playground/src/Core.scala 38:30]
  wire [1:0] Tlb_io_dcache_access_type; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_vpn_ready; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_vpn_valid; // @[playground/src/Core.scala 38:30]
  wire [26:0] Tlb_io_dcache_ptw_vpn_bits; // @[playground/src/Core.scala 38:30]
  wire [1:0] Tlb_io_dcache_ptw_access_type; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_valid; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_page_fault; // @[playground/src/Core.scala 38:30]
  wire [19:0] Tlb_io_dcache_ptw_pte_bits_entry_ppn; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_d; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_g; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_u; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_x; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_w; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_r; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_dcache_ptw_pte_bits_entry_flag_v; // @[playground/src/Core.scala 38:30]
  wire [17:0] Tlb_io_dcache_ptw_pte_bits_rmask; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_dcache_csr_satp; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_dcache_csr_mstatus; // @[playground/src/Core.scala 38:30]
  wire [1:0] Tlb_io_dcache_csr_imode; // @[playground/src/Core.scala 38:30]
  wire [1:0] Tlb_io_dcache_csr_dmode; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_csr_satp; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_csr_mstatus; // @[playground/src/Core.scala 38:30]
  wire [1:0] Tlb_io_csr_imode; // @[playground/src/Core.scala 38:30]
  wire [1:0] Tlb_io_csr_dmode; // @[playground/src/Core.scala 38:30]
  wire  Tlb_io_sfence_vma_valid; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_sfence_vma_src_info_src1_data; // @[playground/src/Core.scala 38:30]
  wire [63:0] Tlb_io_sfence_vma_src_info_src2_data; // @[playground/src/Core.scala 38:30]
  wire [64:0] _T = {{1'd0}, io_inst_addr_0}; // @[playground/src/Core.scala 72:58]
  wire  _T_6 = ~DecodeUnit_io_instFifo_allow_to_go_0 & Ctrl_io_executeUnit_allow_to_go; // @[playground/src/Core.scala 92:43]
  wire  _T_10 = ~DecodeUnit_io_instFifo_allow_to_go_1 & Ctrl_io_executeUnit_allow_to_go; // @[playground/src/Core.scala 92:43]
  Ctrl Ctrl ( // @[playground/src/Core.scala 25:30]
    .io_cacheCtrl_iCache_stall(Ctrl_io_cacheCtrl_iCache_stall),
    .io_fetchUnit_allow_to_go(Ctrl_io_fetchUnit_allow_to_go),
    .io_decodeUnit_inst0_src1_ren(Ctrl_io_decodeUnit_inst0_src1_ren),
    .io_decodeUnit_inst0_src1_raddr(Ctrl_io_decodeUnit_inst0_src1_raddr),
    .io_decodeUnit_inst0_src2_ren(Ctrl_io_decodeUnit_inst0_src2_ren),
    .io_decodeUnit_inst0_src2_raddr(Ctrl_io_decodeUnit_inst0_src2_raddr),
    .io_decodeUnit_branch(Ctrl_io_decodeUnit_branch),
    .io_decodeUnit_allow_to_go(Ctrl_io_decodeUnit_allow_to_go),
    .io_decodeUnit_do_flush(Ctrl_io_decodeUnit_do_flush),
    .io_executeUnit_inst_0_is_load(Ctrl_io_executeUnit_inst_0_is_load),
    .io_executeUnit_inst_0_reg_waddr(Ctrl_io_executeUnit_inst_0_reg_waddr),
    .io_executeUnit_inst_1_is_load(Ctrl_io_executeUnit_inst_1_is_load),
    .io_executeUnit_inst_1_reg_waddr(Ctrl_io_executeUnit_inst_1_reg_waddr),
    .io_executeUnit_flush(Ctrl_io_executeUnit_flush),
    .io_executeUnit_allow_to_go(Ctrl_io_executeUnit_allow_to_go),
    .io_executeUnit_do_flush(Ctrl_io_executeUnit_do_flush),
    .io_executeUnit_fu_allow_to_go(Ctrl_io_executeUnit_fu_allow_to_go),
    .io_executeUnit_fu_stall(Ctrl_io_executeUnit_fu_stall),
    .io_memoryUnit_flush(Ctrl_io_memoryUnit_flush),
    .io_memoryUnit_mem_stall(Ctrl_io_memoryUnit_mem_stall),
    .io_memoryUnit_allow_to_go(Ctrl_io_memoryUnit_allow_to_go),
    .io_memoryUnit_do_flush(Ctrl_io_memoryUnit_do_flush),
    .io_memoryUnit_complete_single_request(Ctrl_io_memoryUnit_complete_single_request),
    .io_writeBackUnit_allow_to_go(Ctrl_io_writeBackUnit_allow_to_go)
  );
  FetchUnit FetchUnit ( // @[playground/src/Core.scala 26:30]
    .clock(FetchUnit_clock),
    .reset(FetchUnit_reset),
    .io_memory_flush(FetchUnit_io_memory_flush),
    .io_memory_target(FetchUnit_io_memory_target),
    .io_decode_branch(FetchUnit_io_decode_branch),
    .io_decode_target(FetchUnit_io_decode_target),
    .io_execute_flush(FetchUnit_io_execute_flush),
    .io_execute_target(FetchUnit_io_execute_target),
    .io_instFifo_full(FetchUnit_io_instFifo_full),
    .io_iCache_inst_valid_0(FetchUnit_io_iCache_inst_valid_0),
    .io_iCache_inst_valid_1(FetchUnit_io_iCache_inst_valid_1),
    .io_iCache_pc(FetchUnit_io_iCache_pc),
    .io_iCache_pc_next(FetchUnit_io_iCache_pc_next)
  );
  BranchPredictorUnit BranchPredictorUnit ( // @[playground/src/Core.scala 27:30]
    .clock(BranchPredictorUnit_clock),
    .reset(BranchPredictorUnit_reset),
    .io_decode_pc(BranchPredictorUnit_io_decode_pc),
    .io_decode_info_valid(BranchPredictorUnit_io_decode_info_valid),
    .io_decode_info_fusel(BranchPredictorUnit_io_decode_info_fusel),
    .io_decode_info_op(BranchPredictorUnit_io_decode_info_op),
    .io_decode_info_imm(BranchPredictorUnit_io_decode_info_imm),
    .io_decode_pht_index(BranchPredictorUnit_io_decode_pht_index),
    .io_decode_branch_inst(BranchPredictorUnit_io_decode_branch_inst),
    .io_decode_branch(BranchPredictorUnit_io_decode_branch),
    .io_decode_target(BranchPredictorUnit_io_decode_target),
    .io_decode_update_pht_index(BranchPredictorUnit_io_decode_update_pht_index),
    .io_instBuffer_pc_0(BranchPredictorUnit_io_instBuffer_pc_0),
    .io_instBuffer_pc_1(BranchPredictorUnit_io_instBuffer_pc_1),
    .io_instBuffer_pht_index_0(BranchPredictorUnit_io_instBuffer_pht_index_0),
    .io_instBuffer_pht_index_1(BranchPredictorUnit_io_instBuffer_pht_index_1),
    .io_execute_pc(BranchPredictorUnit_io_execute_pc),
    .io_execute_update_pht_index(BranchPredictorUnit_io_execute_update_pht_index),
    .io_execute_branch_inst(BranchPredictorUnit_io_execute_branch_inst),
    .io_execute_branch(BranchPredictorUnit_io_execute_branch)
  );
  InstFifo InstFifo ( // @[playground/src/Core.scala 28:30]
    .clock(InstFifo_clock),
    .reset(InstFifo_reset),
    .io_do_flush(InstFifo_io_do_flush),
    .io_wen_0(InstFifo_io_wen_0),
    .io_wen_1(InstFifo_io_wen_1),
    .io_write_0_inst(InstFifo_io_write_0_inst),
    .io_write_0_pht_index(InstFifo_io_write_0_pht_index),
    .io_write_0_addr_misaligned(InstFifo_io_write_0_addr_misaligned),
    .io_write_0_access_fault(InstFifo_io_write_0_access_fault),
    .io_write_0_page_fault(InstFifo_io_write_0_page_fault),
    .io_write_0_pc(InstFifo_io_write_0_pc),
    .io_write_1_inst(InstFifo_io_write_1_inst),
    .io_write_1_pht_index(InstFifo_io_write_1_pht_index),
    .io_write_1_addr_misaligned(InstFifo_io_write_1_addr_misaligned),
    .io_write_1_access_fault(InstFifo_io_write_1_access_fault),
    .io_write_1_page_fault(InstFifo_io_write_1_page_fault),
    .io_write_1_pc(InstFifo_io_write_1_pc),
    .io_full(InstFifo_io_full),
    .io_decoderUint_allow_to_go_0(InstFifo_io_decoderUint_allow_to_go_0),
    .io_decoderUint_allow_to_go_1(InstFifo_io_decoderUint_allow_to_go_1),
    .io_decoderUint_inst_0_inst(InstFifo_io_decoderUint_inst_0_inst),
    .io_decoderUint_inst_0_pht_index(InstFifo_io_decoderUint_inst_0_pht_index),
    .io_decoderUint_inst_0_addr_misaligned(InstFifo_io_decoderUint_inst_0_addr_misaligned),
    .io_decoderUint_inst_0_access_fault(InstFifo_io_decoderUint_inst_0_access_fault),
    .io_decoderUint_inst_0_page_fault(InstFifo_io_decoderUint_inst_0_page_fault),
    .io_decoderUint_inst_0_pc(InstFifo_io_decoderUint_inst_0_pc),
    .io_decoderUint_inst_1_inst(InstFifo_io_decoderUint_inst_1_inst),
    .io_decoderUint_inst_1_addr_misaligned(InstFifo_io_decoderUint_inst_1_addr_misaligned),
    .io_decoderUint_inst_1_access_fault(InstFifo_io_decoderUint_inst_1_access_fault),
    .io_decoderUint_inst_1_page_fault(InstFifo_io_decoderUint_inst_1_page_fault),
    .io_decoderUint_inst_1_pc(InstFifo_io_decoderUint_inst_1_pc),
    .io_decoderUint_info_empty(InstFifo_io_decoderUint_info_empty),
    .io_decoderUint_info_almost_empty(InstFifo_io_decoderUint_info_almost_empty)
  );
  DecodeUnit DecodeUnit ( // @[playground/src/Core.scala 29:30]
    .io_instFifo_allow_to_go_0(DecodeUnit_io_instFifo_allow_to_go_0),
    .io_instFifo_allow_to_go_1(DecodeUnit_io_instFifo_allow_to_go_1),
    .io_instFifo_inst_0_inst(DecodeUnit_io_instFifo_inst_0_inst),
    .io_instFifo_inst_0_pht_index(DecodeUnit_io_instFifo_inst_0_pht_index),
    .io_instFifo_inst_0_addr_misaligned(DecodeUnit_io_instFifo_inst_0_addr_misaligned),
    .io_instFifo_inst_0_access_fault(DecodeUnit_io_instFifo_inst_0_access_fault),
    .io_instFifo_inst_0_page_fault(DecodeUnit_io_instFifo_inst_0_page_fault),
    .io_instFifo_inst_0_pc(DecodeUnit_io_instFifo_inst_0_pc),
    .io_instFifo_inst_1_inst(DecodeUnit_io_instFifo_inst_1_inst),
    .io_instFifo_inst_1_addr_misaligned(DecodeUnit_io_instFifo_inst_1_addr_misaligned),
    .io_instFifo_inst_1_access_fault(DecodeUnit_io_instFifo_inst_1_access_fault),
    .io_instFifo_inst_1_page_fault(DecodeUnit_io_instFifo_inst_1_page_fault),
    .io_instFifo_inst_1_pc(DecodeUnit_io_instFifo_inst_1_pc),
    .io_instFifo_info_empty(DecodeUnit_io_instFifo_info_empty),
    .io_instFifo_info_almost_empty(DecodeUnit_io_instFifo_info_almost_empty),
    .io_regfile_0_src1_raddr(DecodeUnit_io_regfile_0_src1_raddr),
    .io_regfile_0_src1_rdata(DecodeUnit_io_regfile_0_src1_rdata),
    .io_regfile_0_src2_raddr(DecodeUnit_io_regfile_0_src2_raddr),
    .io_regfile_0_src2_rdata(DecodeUnit_io_regfile_0_src2_rdata),
    .io_regfile_1_src1_raddr(DecodeUnit_io_regfile_1_src1_raddr),
    .io_regfile_1_src1_rdata(DecodeUnit_io_regfile_1_src1_rdata),
    .io_regfile_1_src2_raddr(DecodeUnit_io_regfile_1_src2_raddr),
    .io_regfile_1_src2_rdata(DecodeUnit_io_regfile_1_src2_rdata),
    .io_forward_0_exe_wen(DecodeUnit_io_forward_0_exe_wen),
    .io_forward_0_exe_waddr(DecodeUnit_io_forward_0_exe_waddr),
    .io_forward_0_exe_wdata(DecodeUnit_io_forward_0_exe_wdata),
    .io_forward_0_is_load(DecodeUnit_io_forward_0_is_load),
    .io_forward_0_mem_wen(DecodeUnit_io_forward_0_mem_wen),
    .io_forward_0_mem_waddr(DecodeUnit_io_forward_0_mem_waddr),
    .io_forward_0_mem_wdata(DecodeUnit_io_forward_0_mem_wdata),
    .io_forward_1_exe_wen(DecodeUnit_io_forward_1_exe_wen),
    .io_forward_1_exe_waddr(DecodeUnit_io_forward_1_exe_waddr),
    .io_forward_1_exe_wdata(DecodeUnit_io_forward_1_exe_wdata),
    .io_forward_1_is_load(DecodeUnit_io_forward_1_is_load),
    .io_forward_1_mem_wen(DecodeUnit_io_forward_1_mem_wen),
    .io_forward_1_mem_waddr(DecodeUnit_io_forward_1_mem_waddr),
    .io_forward_1_mem_wdata(DecodeUnit_io_forward_1_mem_wdata),
    .io_csr_mode(DecodeUnit_io_csr_mode),
    .io_csr_interrupt(DecodeUnit_io_csr_interrupt),
    .io_fetchUnit_branch(DecodeUnit_io_fetchUnit_branch),
    .io_fetchUnit_target(DecodeUnit_io_fetchUnit_target),
    .io_bpu_pc(DecodeUnit_io_bpu_pc),
    .io_bpu_info_valid(DecodeUnit_io_bpu_info_valid),
    .io_bpu_info_fusel(DecodeUnit_io_bpu_info_fusel),
    .io_bpu_info_op(DecodeUnit_io_bpu_info_op),
    .io_bpu_info_imm(DecodeUnit_io_bpu_info_imm),
    .io_bpu_pht_index(DecodeUnit_io_bpu_pht_index),
    .io_bpu_branch_inst(DecodeUnit_io_bpu_branch_inst),
    .io_bpu_branch(DecodeUnit_io_bpu_branch),
    .io_bpu_target(DecodeUnit_io_bpu_target),
    .io_bpu_update_pht_index(DecodeUnit_io_bpu_update_pht_index),
    .io_executeStage_inst_0_pc(DecodeUnit_io_executeStage_inst_0_pc),
    .io_executeStage_inst_0_info_valid(DecodeUnit_io_executeStage_inst_0_info_valid),
    .io_executeStage_inst_0_info_fusel(DecodeUnit_io_executeStage_inst_0_info_fusel),
    .io_executeStage_inst_0_info_op(DecodeUnit_io_executeStage_inst_0_info_op),
    .io_executeStage_inst_0_info_reg_wen(DecodeUnit_io_executeStage_inst_0_info_reg_wen),
    .io_executeStage_inst_0_info_reg_waddr(DecodeUnit_io_executeStage_inst_0_info_reg_waddr),
    .io_executeStage_inst_0_info_imm(DecodeUnit_io_executeStage_inst_0_info_imm),
    .io_executeStage_inst_0_info_inst(DecodeUnit_io_executeStage_inst_0_info_inst),
    .io_executeStage_inst_0_src_info_src1_data(DecodeUnit_io_executeStage_inst_0_src_info_src1_data),
    .io_executeStage_inst_0_src_info_src2_data(DecodeUnit_io_executeStage_inst_0_src_info_src2_data),
    .io_executeStage_inst_0_ex_exception_0(DecodeUnit_io_executeStage_inst_0_ex_exception_0),
    .io_executeStage_inst_0_ex_exception_1(DecodeUnit_io_executeStage_inst_0_ex_exception_1),
    .io_executeStage_inst_0_ex_exception_2(DecodeUnit_io_executeStage_inst_0_ex_exception_2),
    .io_executeStage_inst_0_ex_exception_3(DecodeUnit_io_executeStage_inst_0_ex_exception_3),
    .io_executeStage_inst_0_ex_exception_8(DecodeUnit_io_executeStage_inst_0_ex_exception_8),
    .io_executeStage_inst_0_ex_exception_9(DecodeUnit_io_executeStage_inst_0_ex_exception_9),
    .io_executeStage_inst_0_ex_exception_11(DecodeUnit_io_executeStage_inst_0_ex_exception_11),
    .io_executeStage_inst_0_ex_exception_12(DecodeUnit_io_executeStage_inst_0_ex_exception_12),
    .io_executeStage_inst_0_ex_interrupt_0(DecodeUnit_io_executeStage_inst_0_ex_interrupt_0),
    .io_executeStage_inst_0_ex_interrupt_1(DecodeUnit_io_executeStage_inst_0_ex_interrupt_1),
    .io_executeStage_inst_0_ex_interrupt_2(DecodeUnit_io_executeStage_inst_0_ex_interrupt_2),
    .io_executeStage_inst_0_ex_interrupt_3(DecodeUnit_io_executeStage_inst_0_ex_interrupt_3),
    .io_executeStage_inst_0_ex_interrupt_4(DecodeUnit_io_executeStage_inst_0_ex_interrupt_4),
    .io_executeStage_inst_0_ex_interrupt_5(DecodeUnit_io_executeStage_inst_0_ex_interrupt_5),
    .io_executeStage_inst_0_ex_interrupt_6(DecodeUnit_io_executeStage_inst_0_ex_interrupt_6),
    .io_executeStage_inst_0_ex_interrupt_7(DecodeUnit_io_executeStage_inst_0_ex_interrupt_7),
    .io_executeStage_inst_0_ex_interrupt_8(DecodeUnit_io_executeStage_inst_0_ex_interrupt_8),
    .io_executeStage_inst_0_ex_interrupt_9(DecodeUnit_io_executeStage_inst_0_ex_interrupt_9),
    .io_executeStage_inst_0_ex_interrupt_10(DecodeUnit_io_executeStage_inst_0_ex_interrupt_10),
    .io_executeStage_inst_0_ex_interrupt_11(DecodeUnit_io_executeStage_inst_0_ex_interrupt_11),
    .io_executeStage_inst_0_ex_tval_0(DecodeUnit_io_executeStage_inst_0_ex_tval_0),
    .io_executeStage_inst_0_ex_tval_1(DecodeUnit_io_executeStage_inst_0_ex_tval_1),
    .io_executeStage_inst_0_ex_tval_2(DecodeUnit_io_executeStage_inst_0_ex_tval_2),
    .io_executeStage_inst_0_ex_tval_12(DecodeUnit_io_executeStage_inst_0_ex_tval_12),
    .io_executeStage_inst_1_pc(DecodeUnit_io_executeStage_inst_1_pc),
    .io_executeStage_inst_1_info_valid(DecodeUnit_io_executeStage_inst_1_info_valid),
    .io_executeStage_inst_1_info_fusel(DecodeUnit_io_executeStage_inst_1_info_fusel),
    .io_executeStage_inst_1_info_op(DecodeUnit_io_executeStage_inst_1_info_op),
    .io_executeStage_inst_1_info_reg_wen(DecodeUnit_io_executeStage_inst_1_info_reg_wen),
    .io_executeStage_inst_1_info_reg_waddr(DecodeUnit_io_executeStage_inst_1_info_reg_waddr),
    .io_executeStage_inst_1_info_imm(DecodeUnit_io_executeStage_inst_1_info_imm),
    .io_executeStage_inst_1_info_inst(DecodeUnit_io_executeStage_inst_1_info_inst),
    .io_executeStage_inst_1_src_info_src1_data(DecodeUnit_io_executeStage_inst_1_src_info_src1_data),
    .io_executeStage_inst_1_src_info_src2_data(DecodeUnit_io_executeStage_inst_1_src_info_src2_data),
    .io_executeStage_inst_1_ex_exception_0(DecodeUnit_io_executeStage_inst_1_ex_exception_0),
    .io_executeStage_inst_1_ex_exception_1(DecodeUnit_io_executeStage_inst_1_ex_exception_1),
    .io_executeStage_inst_1_ex_exception_2(DecodeUnit_io_executeStage_inst_1_ex_exception_2),
    .io_executeStage_inst_1_ex_exception_3(DecodeUnit_io_executeStage_inst_1_ex_exception_3),
    .io_executeStage_inst_1_ex_exception_8(DecodeUnit_io_executeStage_inst_1_ex_exception_8),
    .io_executeStage_inst_1_ex_exception_9(DecodeUnit_io_executeStage_inst_1_ex_exception_9),
    .io_executeStage_inst_1_ex_exception_11(DecodeUnit_io_executeStage_inst_1_ex_exception_11),
    .io_executeStage_inst_1_ex_exception_12(DecodeUnit_io_executeStage_inst_1_ex_exception_12),
    .io_executeStage_inst_1_ex_interrupt_0(DecodeUnit_io_executeStage_inst_1_ex_interrupt_0),
    .io_executeStage_inst_1_ex_interrupt_1(DecodeUnit_io_executeStage_inst_1_ex_interrupt_1),
    .io_executeStage_inst_1_ex_interrupt_2(DecodeUnit_io_executeStage_inst_1_ex_interrupt_2),
    .io_executeStage_inst_1_ex_interrupt_3(DecodeUnit_io_executeStage_inst_1_ex_interrupt_3),
    .io_executeStage_inst_1_ex_interrupt_4(DecodeUnit_io_executeStage_inst_1_ex_interrupt_4),
    .io_executeStage_inst_1_ex_interrupt_5(DecodeUnit_io_executeStage_inst_1_ex_interrupt_5),
    .io_executeStage_inst_1_ex_interrupt_6(DecodeUnit_io_executeStage_inst_1_ex_interrupt_6),
    .io_executeStage_inst_1_ex_interrupt_7(DecodeUnit_io_executeStage_inst_1_ex_interrupt_7),
    .io_executeStage_inst_1_ex_interrupt_8(DecodeUnit_io_executeStage_inst_1_ex_interrupt_8),
    .io_executeStage_inst_1_ex_interrupt_9(DecodeUnit_io_executeStage_inst_1_ex_interrupt_9),
    .io_executeStage_inst_1_ex_interrupt_10(DecodeUnit_io_executeStage_inst_1_ex_interrupt_10),
    .io_executeStage_inst_1_ex_interrupt_11(DecodeUnit_io_executeStage_inst_1_ex_interrupt_11),
    .io_executeStage_inst_1_ex_tval_0(DecodeUnit_io_executeStage_inst_1_ex_tval_0),
    .io_executeStage_inst_1_ex_tval_1(DecodeUnit_io_executeStage_inst_1_ex_tval_1),
    .io_executeStage_inst_1_ex_tval_2(DecodeUnit_io_executeStage_inst_1_ex_tval_2),
    .io_executeStage_inst_1_ex_tval_12(DecodeUnit_io_executeStage_inst_1_ex_tval_12),
    .io_executeStage_jump_branch_info_jump_regiser(DecodeUnit_io_executeStage_jump_branch_info_jump_regiser),
    .io_executeStage_jump_branch_info_branch_inst(DecodeUnit_io_executeStage_jump_branch_info_branch_inst),
    .io_executeStage_jump_branch_info_pred_branch(DecodeUnit_io_executeStage_jump_branch_info_pred_branch),
    .io_executeStage_jump_branch_info_branch_target(DecodeUnit_io_executeStage_jump_branch_info_branch_target),
    .io_executeStage_jump_branch_info_update_pht_index(DecodeUnit_io_executeStage_jump_branch_info_update_pht_index),
    .io_ctrl_inst0_src1_ren(DecodeUnit_io_ctrl_inst0_src1_ren),
    .io_ctrl_inst0_src1_raddr(DecodeUnit_io_ctrl_inst0_src1_raddr),
    .io_ctrl_inst0_src2_ren(DecodeUnit_io_ctrl_inst0_src2_ren),
    .io_ctrl_inst0_src2_raddr(DecodeUnit_io_ctrl_inst0_src2_raddr),
    .io_ctrl_branch(DecodeUnit_io_ctrl_branch),
    .io_ctrl_allow_to_go(DecodeUnit_io_ctrl_allow_to_go)
  );
  ARegFile ARegFile ( // @[playground/src/Core.scala 30:30]
    .clock(ARegFile_clock),
    .reset(ARegFile_reset),
    .io_read_0_src1_raddr(ARegFile_io_read_0_src1_raddr),
    .io_read_0_src1_rdata(ARegFile_io_read_0_src1_rdata),
    .io_read_0_src2_raddr(ARegFile_io_read_0_src2_raddr),
    .io_read_0_src2_rdata(ARegFile_io_read_0_src2_rdata),
    .io_read_1_src1_raddr(ARegFile_io_read_1_src1_raddr),
    .io_read_1_src1_rdata(ARegFile_io_read_1_src1_rdata),
    .io_read_1_src2_raddr(ARegFile_io_read_1_src2_raddr),
    .io_read_1_src2_rdata(ARegFile_io_read_1_src2_rdata),
    .io_write_0_wen(ARegFile_io_write_0_wen),
    .io_write_0_waddr(ARegFile_io_write_0_waddr),
    .io_write_0_wdata(ARegFile_io_write_0_wdata),
    .io_write_1_wen(ARegFile_io_write_1_wen),
    .io_write_1_waddr(ARegFile_io_write_1_waddr),
    .io_write_1_wdata(ARegFile_io_write_1_wdata)
  );
  ExecuteStage ExecuteStage ( // @[playground/src/Core.scala 31:30]
    .clock(ExecuteStage_clock),
    .reset(ExecuteStage_reset),
    .io_ctrl_allow_to_go_0(ExecuteStage_io_ctrl_allow_to_go_0),
    .io_ctrl_allow_to_go_1(ExecuteStage_io_ctrl_allow_to_go_1),
    .io_ctrl_clear_0(ExecuteStage_io_ctrl_clear_0),
    .io_ctrl_clear_1(ExecuteStage_io_ctrl_clear_1),
    .io_decodeUnit_inst_0_pc(ExecuteStage_io_decodeUnit_inst_0_pc),
    .io_decodeUnit_inst_0_info_valid(ExecuteStage_io_decodeUnit_inst_0_info_valid),
    .io_decodeUnit_inst_0_info_fusel(ExecuteStage_io_decodeUnit_inst_0_info_fusel),
    .io_decodeUnit_inst_0_info_op(ExecuteStage_io_decodeUnit_inst_0_info_op),
    .io_decodeUnit_inst_0_info_reg_wen(ExecuteStage_io_decodeUnit_inst_0_info_reg_wen),
    .io_decodeUnit_inst_0_info_reg_waddr(ExecuteStage_io_decodeUnit_inst_0_info_reg_waddr),
    .io_decodeUnit_inst_0_info_imm(ExecuteStage_io_decodeUnit_inst_0_info_imm),
    .io_decodeUnit_inst_0_info_inst(ExecuteStage_io_decodeUnit_inst_0_info_inst),
    .io_decodeUnit_inst_0_src_info_src1_data(ExecuteStage_io_decodeUnit_inst_0_src_info_src1_data),
    .io_decodeUnit_inst_0_src_info_src2_data(ExecuteStage_io_decodeUnit_inst_0_src_info_src2_data),
    .io_decodeUnit_inst_0_ex_exception_0(ExecuteStage_io_decodeUnit_inst_0_ex_exception_0),
    .io_decodeUnit_inst_0_ex_exception_1(ExecuteStage_io_decodeUnit_inst_0_ex_exception_1),
    .io_decodeUnit_inst_0_ex_exception_2(ExecuteStage_io_decodeUnit_inst_0_ex_exception_2),
    .io_decodeUnit_inst_0_ex_exception_3(ExecuteStage_io_decodeUnit_inst_0_ex_exception_3),
    .io_decodeUnit_inst_0_ex_exception_8(ExecuteStage_io_decodeUnit_inst_0_ex_exception_8),
    .io_decodeUnit_inst_0_ex_exception_9(ExecuteStage_io_decodeUnit_inst_0_ex_exception_9),
    .io_decodeUnit_inst_0_ex_exception_11(ExecuteStage_io_decodeUnit_inst_0_ex_exception_11),
    .io_decodeUnit_inst_0_ex_exception_12(ExecuteStage_io_decodeUnit_inst_0_ex_exception_12),
    .io_decodeUnit_inst_0_ex_interrupt_0(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_0),
    .io_decodeUnit_inst_0_ex_interrupt_1(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_1),
    .io_decodeUnit_inst_0_ex_interrupt_2(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_2),
    .io_decodeUnit_inst_0_ex_interrupt_3(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_3),
    .io_decodeUnit_inst_0_ex_interrupt_4(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_4),
    .io_decodeUnit_inst_0_ex_interrupt_5(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_5),
    .io_decodeUnit_inst_0_ex_interrupt_6(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_6),
    .io_decodeUnit_inst_0_ex_interrupt_7(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_7),
    .io_decodeUnit_inst_0_ex_interrupt_8(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_8),
    .io_decodeUnit_inst_0_ex_interrupt_9(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_9),
    .io_decodeUnit_inst_0_ex_interrupt_10(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_10),
    .io_decodeUnit_inst_0_ex_interrupt_11(ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_11),
    .io_decodeUnit_inst_0_ex_tval_0(ExecuteStage_io_decodeUnit_inst_0_ex_tval_0),
    .io_decodeUnit_inst_0_ex_tval_1(ExecuteStage_io_decodeUnit_inst_0_ex_tval_1),
    .io_decodeUnit_inst_0_ex_tval_2(ExecuteStage_io_decodeUnit_inst_0_ex_tval_2),
    .io_decodeUnit_inst_0_ex_tval_12(ExecuteStage_io_decodeUnit_inst_0_ex_tval_12),
    .io_decodeUnit_inst_1_pc(ExecuteStage_io_decodeUnit_inst_1_pc),
    .io_decodeUnit_inst_1_info_valid(ExecuteStage_io_decodeUnit_inst_1_info_valid),
    .io_decodeUnit_inst_1_info_fusel(ExecuteStage_io_decodeUnit_inst_1_info_fusel),
    .io_decodeUnit_inst_1_info_op(ExecuteStage_io_decodeUnit_inst_1_info_op),
    .io_decodeUnit_inst_1_info_reg_wen(ExecuteStage_io_decodeUnit_inst_1_info_reg_wen),
    .io_decodeUnit_inst_1_info_reg_waddr(ExecuteStage_io_decodeUnit_inst_1_info_reg_waddr),
    .io_decodeUnit_inst_1_info_imm(ExecuteStage_io_decodeUnit_inst_1_info_imm),
    .io_decodeUnit_inst_1_info_inst(ExecuteStage_io_decodeUnit_inst_1_info_inst),
    .io_decodeUnit_inst_1_src_info_src1_data(ExecuteStage_io_decodeUnit_inst_1_src_info_src1_data),
    .io_decodeUnit_inst_1_src_info_src2_data(ExecuteStage_io_decodeUnit_inst_1_src_info_src2_data),
    .io_decodeUnit_inst_1_ex_exception_0(ExecuteStage_io_decodeUnit_inst_1_ex_exception_0),
    .io_decodeUnit_inst_1_ex_exception_1(ExecuteStage_io_decodeUnit_inst_1_ex_exception_1),
    .io_decodeUnit_inst_1_ex_exception_2(ExecuteStage_io_decodeUnit_inst_1_ex_exception_2),
    .io_decodeUnit_inst_1_ex_exception_3(ExecuteStage_io_decodeUnit_inst_1_ex_exception_3),
    .io_decodeUnit_inst_1_ex_exception_8(ExecuteStage_io_decodeUnit_inst_1_ex_exception_8),
    .io_decodeUnit_inst_1_ex_exception_9(ExecuteStage_io_decodeUnit_inst_1_ex_exception_9),
    .io_decodeUnit_inst_1_ex_exception_11(ExecuteStage_io_decodeUnit_inst_1_ex_exception_11),
    .io_decodeUnit_inst_1_ex_exception_12(ExecuteStage_io_decodeUnit_inst_1_ex_exception_12),
    .io_decodeUnit_inst_1_ex_interrupt_0(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_0),
    .io_decodeUnit_inst_1_ex_interrupt_1(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_1),
    .io_decodeUnit_inst_1_ex_interrupt_2(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_2),
    .io_decodeUnit_inst_1_ex_interrupt_3(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_3),
    .io_decodeUnit_inst_1_ex_interrupt_4(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_4),
    .io_decodeUnit_inst_1_ex_interrupt_5(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_5),
    .io_decodeUnit_inst_1_ex_interrupt_6(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_6),
    .io_decodeUnit_inst_1_ex_interrupt_7(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_7),
    .io_decodeUnit_inst_1_ex_interrupt_8(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_8),
    .io_decodeUnit_inst_1_ex_interrupt_9(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_9),
    .io_decodeUnit_inst_1_ex_interrupt_10(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_10),
    .io_decodeUnit_inst_1_ex_interrupt_11(ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_11),
    .io_decodeUnit_inst_1_ex_tval_0(ExecuteStage_io_decodeUnit_inst_1_ex_tval_0),
    .io_decodeUnit_inst_1_ex_tval_1(ExecuteStage_io_decodeUnit_inst_1_ex_tval_1),
    .io_decodeUnit_inst_1_ex_tval_2(ExecuteStage_io_decodeUnit_inst_1_ex_tval_2),
    .io_decodeUnit_inst_1_ex_tval_12(ExecuteStage_io_decodeUnit_inst_1_ex_tval_12),
    .io_decodeUnit_jump_branch_info_jump_regiser(ExecuteStage_io_decodeUnit_jump_branch_info_jump_regiser),
    .io_decodeUnit_jump_branch_info_branch_inst(ExecuteStage_io_decodeUnit_jump_branch_info_branch_inst),
    .io_decodeUnit_jump_branch_info_pred_branch(ExecuteStage_io_decodeUnit_jump_branch_info_pred_branch),
    .io_decodeUnit_jump_branch_info_branch_target(ExecuteStage_io_decodeUnit_jump_branch_info_branch_target),
    .io_decodeUnit_jump_branch_info_update_pht_index(ExecuteStage_io_decodeUnit_jump_branch_info_update_pht_index),
    .io_executeUnit_inst_0_pc(ExecuteStage_io_executeUnit_inst_0_pc),
    .io_executeUnit_inst_0_info_valid(ExecuteStage_io_executeUnit_inst_0_info_valid),
    .io_executeUnit_inst_0_info_fusel(ExecuteStage_io_executeUnit_inst_0_info_fusel),
    .io_executeUnit_inst_0_info_op(ExecuteStage_io_executeUnit_inst_0_info_op),
    .io_executeUnit_inst_0_info_reg_wen(ExecuteStage_io_executeUnit_inst_0_info_reg_wen),
    .io_executeUnit_inst_0_info_reg_waddr(ExecuteStage_io_executeUnit_inst_0_info_reg_waddr),
    .io_executeUnit_inst_0_info_imm(ExecuteStage_io_executeUnit_inst_0_info_imm),
    .io_executeUnit_inst_0_info_inst(ExecuteStage_io_executeUnit_inst_0_info_inst),
    .io_executeUnit_inst_0_src_info_src1_data(ExecuteStage_io_executeUnit_inst_0_src_info_src1_data),
    .io_executeUnit_inst_0_src_info_src2_data(ExecuteStage_io_executeUnit_inst_0_src_info_src2_data),
    .io_executeUnit_inst_0_ex_exception_0(ExecuteStage_io_executeUnit_inst_0_ex_exception_0),
    .io_executeUnit_inst_0_ex_exception_1(ExecuteStage_io_executeUnit_inst_0_ex_exception_1),
    .io_executeUnit_inst_0_ex_exception_2(ExecuteStage_io_executeUnit_inst_0_ex_exception_2),
    .io_executeUnit_inst_0_ex_exception_3(ExecuteStage_io_executeUnit_inst_0_ex_exception_3),
    .io_executeUnit_inst_0_ex_exception_8(ExecuteStage_io_executeUnit_inst_0_ex_exception_8),
    .io_executeUnit_inst_0_ex_exception_9(ExecuteStage_io_executeUnit_inst_0_ex_exception_9),
    .io_executeUnit_inst_0_ex_exception_11(ExecuteStage_io_executeUnit_inst_0_ex_exception_11),
    .io_executeUnit_inst_0_ex_exception_12(ExecuteStage_io_executeUnit_inst_0_ex_exception_12),
    .io_executeUnit_inst_0_ex_interrupt_0(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_0),
    .io_executeUnit_inst_0_ex_interrupt_1(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_1),
    .io_executeUnit_inst_0_ex_interrupt_2(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_2),
    .io_executeUnit_inst_0_ex_interrupt_3(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_3),
    .io_executeUnit_inst_0_ex_interrupt_4(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_4),
    .io_executeUnit_inst_0_ex_interrupt_5(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_5),
    .io_executeUnit_inst_0_ex_interrupt_6(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_6),
    .io_executeUnit_inst_0_ex_interrupt_7(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_7),
    .io_executeUnit_inst_0_ex_interrupt_8(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_8),
    .io_executeUnit_inst_0_ex_interrupt_9(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_9),
    .io_executeUnit_inst_0_ex_interrupt_10(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_10),
    .io_executeUnit_inst_0_ex_interrupt_11(ExecuteStage_io_executeUnit_inst_0_ex_interrupt_11),
    .io_executeUnit_inst_0_ex_tval_0(ExecuteStage_io_executeUnit_inst_0_ex_tval_0),
    .io_executeUnit_inst_0_ex_tval_1(ExecuteStage_io_executeUnit_inst_0_ex_tval_1),
    .io_executeUnit_inst_0_ex_tval_2(ExecuteStage_io_executeUnit_inst_0_ex_tval_2),
    .io_executeUnit_inst_0_ex_tval_12(ExecuteStage_io_executeUnit_inst_0_ex_tval_12),
    .io_executeUnit_inst_1_pc(ExecuteStage_io_executeUnit_inst_1_pc),
    .io_executeUnit_inst_1_info_valid(ExecuteStage_io_executeUnit_inst_1_info_valid),
    .io_executeUnit_inst_1_info_fusel(ExecuteStage_io_executeUnit_inst_1_info_fusel),
    .io_executeUnit_inst_1_info_op(ExecuteStage_io_executeUnit_inst_1_info_op),
    .io_executeUnit_inst_1_info_reg_wen(ExecuteStage_io_executeUnit_inst_1_info_reg_wen),
    .io_executeUnit_inst_1_info_reg_waddr(ExecuteStage_io_executeUnit_inst_1_info_reg_waddr),
    .io_executeUnit_inst_1_info_imm(ExecuteStage_io_executeUnit_inst_1_info_imm),
    .io_executeUnit_inst_1_info_inst(ExecuteStage_io_executeUnit_inst_1_info_inst),
    .io_executeUnit_inst_1_src_info_src1_data(ExecuteStage_io_executeUnit_inst_1_src_info_src1_data),
    .io_executeUnit_inst_1_src_info_src2_data(ExecuteStage_io_executeUnit_inst_1_src_info_src2_data),
    .io_executeUnit_inst_1_ex_exception_0(ExecuteStage_io_executeUnit_inst_1_ex_exception_0),
    .io_executeUnit_inst_1_ex_exception_1(ExecuteStage_io_executeUnit_inst_1_ex_exception_1),
    .io_executeUnit_inst_1_ex_exception_2(ExecuteStage_io_executeUnit_inst_1_ex_exception_2),
    .io_executeUnit_inst_1_ex_exception_3(ExecuteStage_io_executeUnit_inst_1_ex_exception_3),
    .io_executeUnit_inst_1_ex_exception_8(ExecuteStage_io_executeUnit_inst_1_ex_exception_8),
    .io_executeUnit_inst_1_ex_exception_9(ExecuteStage_io_executeUnit_inst_1_ex_exception_9),
    .io_executeUnit_inst_1_ex_exception_11(ExecuteStage_io_executeUnit_inst_1_ex_exception_11),
    .io_executeUnit_inst_1_ex_exception_12(ExecuteStage_io_executeUnit_inst_1_ex_exception_12),
    .io_executeUnit_inst_1_ex_interrupt_0(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_0),
    .io_executeUnit_inst_1_ex_interrupt_1(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_1),
    .io_executeUnit_inst_1_ex_interrupt_2(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_2),
    .io_executeUnit_inst_1_ex_interrupt_3(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_3),
    .io_executeUnit_inst_1_ex_interrupt_4(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_4),
    .io_executeUnit_inst_1_ex_interrupt_5(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_5),
    .io_executeUnit_inst_1_ex_interrupt_6(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_6),
    .io_executeUnit_inst_1_ex_interrupt_7(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_7),
    .io_executeUnit_inst_1_ex_interrupt_8(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_8),
    .io_executeUnit_inst_1_ex_interrupt_9(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_9),
    .io_executeUnit_inst_1_ex_interrupt_10(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_10),
    .io_executeUnit_inst_1_ex_interrupt_11(ExecuteStage_io_executeUnit_inst_1_ex_interrupt_11),
    .io_executeUnit_inst_1_ex_tval_0(ExecuteStage_io_executeUnit_inst_1_ex_tval_0),
    .io_executeUnit_inst_1_ex_tval_1(ExecuteStage_io_executeUnit_inst_1_ex_tval_1),
    .io_executeUnit_inst_1_ex_tval_2(ExecuteStage_io_executeUnit_inst_1_ex_tval_2),
    .io_executeUnit_inst_1_ex_tval_12(ExecuteStage_io_executeUnit_inst_1_ex_tval_12),
    .io_executeUnit_jump_branch_info_jump_regiser(ExecuteStage_io_executeUnit_jump_branch_info_jump_regiser),
    .io_executeUnit_jump_branch_info_branch_inst(ExecuteStage_io_executeUnit_jump_branch_info_branch_inst),
    .io_executeUnit_jump_branch_info_pred_branch(ExecuteStage_io_executeUnit_jump_branch_info_pred_branch),
    .io_executeUnit_jump_branch_info_branch_target(ExecuteStage_io_executeUnit_jump_branch_info_branch_target),
    .io_executeUnit_jump_branch_info_update_pht_index(ExecuteStage_io_executeUnit_jump_branch_info_update_pht_index)
  );
  ExecuteUnit ExecuteUnit ( // @[playground/src/Core.scala 32:30]
    .clock(ExecuteUnit_clock),
    .reset(ExecuteUnit_reset),
    .io_ctrl_inst_0_is_load(ExecuteUnit_io_ctrl_inst_0_is_load),
    .io_ctrl_inst_0_reg_waddr(ExecuteUnit_io_ctrl_inst_0_reg_waddr),
    .io_ctrl_inst_1_is_load(ExecuteUnit_io_ctrl_inst_1_is_load),
    .io_ctrl_inst_1_reg_waddr(ExecuteUnit_io_ctrl_inst_1_reg_waddr),
    .io_ctrl_flush(ExecuteUnit_io_ctrl_flush),
    .io_ctrl_allow_to_go(ExecuteUnit_io_ctrl_allow_to_go),
    .io_ctrl_fu_allow_to_go(ExecuteUnit_io_ctrl_fu_allow_to_go),
    .io_ctrl_fu_stall(ExecuteUnit_io_ctrl_fu_stall),
    .io_executeStage_inst_0_pc(ExecuteUnit_io_executeStage_inst_0_pc),
    .io_executeStage_inst_0_info_valid(ExecuteUnit_io_executeStage_inst_0_info_valid),
    .io_executeStage_inst_0_info_fusel(ExecuteUnit_io_executeStage_inst_0_info_fusel),
    .io_executeStage_inst_0_info_op(ExecuteUnit_io_executeStage_inst_0_info_op),
    .io_executeStage_inst_0_info_reg_wen(ExecuteUnit_io_executeStage_inst_0_info_reg_wen),
    .io_executeStage_inst_0_info_reg_waddr(ExecuteUnit_io_executeStage_inst_0_info_reg_waddr),
    .io_executeStage_inst_0_info_imm(ExecuteUnit_io_executeStage_inst_0_info_imm),
    .io_executeStage_inst_0_info_inst(ExecuteUnit_io_executeStage_inst_0_info_inst),
    .io_executeStage_inst_0_src_info_src1_data(ExecuteUnit_io_executeStage_inst_0_src_info_src1_data),
    .io_executeStage_inst_0_src_info_src2_data(ExecuteUnit_io_executeStage_inst_0_src_info_src2_data),
    .io_executeStage_inst_0_ex_exception_0(ExecuteUnit_io_executeStage_inst_0_ex_exception_0),
    .io_executeStage_inst_0_ex_exception_1(ExecuteUnit_io_executeStage_inst_0_ex_exception_1),
    .io_executeStage_inst_0_ex_exception_2(ExecuteUnit_io_executeStage_inst_0_ex_exception_2),
    .io_executeStage_inst_0_ex_exception_3(ExecuteUnit_io_executeStage_inst_0_ex_exception_3),
    .io_executeStage_inst_0_ex_exception_8(ExecuteUnit_io_executeStage_inst_0_ex_exception_8),
    .io_executeStage_inst_0_ex_exception_9(ExecuteUnit_io_executeStage_inst_0_ex_exception_9),
    .io_executeStage_inst_0_ex_exception_11(ExecuteUnit_io_executeStage_inst_0_ex_exception_11),
    .io_executeStage_inst_0_ex_exception_12(ExecuteUnit_io_executeStage_inst_0_ex_exception_12),
    .io_executeStage_inst_0_ex_interrupt_0(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_0),
    .io_executeStage_inst_0_ex_interrupt_1(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_1),
    .io_executeStage_inst_0_ex_interrupt_2(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_2),
    .io_executeStage_inst_0_ex_interrupt_3(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_3),
    .io_executeStage_inst_0_ex_interrupt_4(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_4),
    .io_executeStage_inst_0_ex_interrupt_5(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_5),
    .io_executeStage_inst_0_ex_interrupt_6(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_6),
    .io_executeStage_inst_0_ex_interrupt_7(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_7),
    .io_executeStage_inst_0_ex_interrupt_8(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_8),
    .io_executeStage_inst_0_ex_interrupt_9(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_9),
    .io_executeStage_inst_0_ex_interrupt_10(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_10),
    .io_executeStage_inst_0_ex_interrupt_11(ExecuteUnit_io_executeStage_inst_0_ex_interrupt_11),
    .io_executeStage_inst_0_ex_tval_0(ExecuteUnit_io_executeStage_inst_0_ex_tval_0),
    .io_executeStage_inst_0_ex_tval_1(ExecuteUnit_io_executeStage_inst_0_ex_tval_1),
    .io_executeStage_inst_0_ex_tval_2(ExecuteUnit_io_executeStage_inst_0_ex_tval_2),
    .io_executeStage_inst_0_ex_tval_12(ExecuteUnit_io_executeStage_inst_0_ex_tval_12),
    .io_executeStage_inst_1_pc(ExecuteUnit_io_executeStage_inst_1_pc),
    .io_executeStage_inst_1_info_valid(ExecuteUnit_io_executeStage_inst_1_info_valid),
    .io_executeStage_inst_1_info_fusel(ExecuteUnit_io_executeStage_inst_1_info_fusel),
    .io_executeStage_inst_1_info_op(ExecuteUnit_io_executeStage_inst_1_info_op),
    .io_executeStage_inst_1_info_reg_wen(ExecuteUnit_io_executeStage_inst_1_info_reg_wen),
    .io_executeStage_inst_1_info_reg_waddr(ExecuteUnit_io_executeStage_inst_1_info_reg_waddr),
    .io_executeStage_inst_1_info_imm(ExecuteUnit_io_executeStage_inst_1_info_imm),
    .io_executeStage_inst_1_info_inst(ExecuteUnit_io_executeStage_inst_1_info_inst),
    .io_executeStage_inst_1_src_info_src1_data(ExecuteUnit_io_executeStage_inst_1_src_info_src1_data),
    .io_executeStage_inst_1_src_info_src2_data(ExecuteUnit_io_executeStage_inst_1_src_info_src2_data),
    .io_executeStage_inst_1_ex_exception_0(ExecuteUnit_io_executeStage_inst_1_ex_exception_0),
    .io_executeStage_inst_1_ex_exception_1(ExecuteUnit_io_executeStage_inst_1_ex_exception_1),
    .io_executeStage_inst_1_ex_exception_2(ExecuteUnit_io_executeStage_inst_1_ex_exception_2),
    .io_executeStage_inst_1_ex_exception_3(ExecuteUnit_io_executeStage_inst_1_ex_exception_3),
    .io_executeStage_inst_1_ex_exception_8(ExecuteUnit_io_executeStage_inst_1_ex_exception_8),
    .io_executeStage_inst_1_ex_exception_9(ExecuteUnit_io_executeStage_inst_1_ex_exception_9),
    .io_executeStage_inst_1_ex_exception_11(ExecuteUnit_io_executeStage_inst_1_ex_exception_11),
    .io_executeStage_inst_1_ex_exception_12(ExecuteUnit_io_executeStage_inst_1_ex_exception_12),
    .io_executeStage_inst_1_ex_interrupt_0(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_0),
    .io_executeStage_inst_1_ex_interrupt_1(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_1),
    .io_executeStage_inst_1_ex_interrupt_2(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_2),
    .io_executeStage_inst_1_ex_interrupt_3(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_3),
    .io_executeStage_inst_1_ex_interrupt_4(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_4),
    .io_executeStage_inst_1_ex_interrupt_5(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_5),
    .io_executeStage_inst_1_ex_interrupt_6(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_6),
    .io_executeStage_inst_1_ex_interrupt_7(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_7),
    .io_executeStage_inst_1_ex_interrupt_8(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_8),
    .io_executeStage_inst_1_ex_interrupt_9(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_9),
    .io_executeStage_inst_1_ex_interrupt_10(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_10),
    .io_executeStage_inst_1_ex_interrupt_11(ExecuteUnit_io_executeStage_inst_1_ex_interrupt_11),
    .io_executeStage_inst_1_ex_tval_0(ExecuteUnit_io_executeStage_inst_1_ex_tval_0),
    .io_executeStage_inst_1_ex_tval_1(ExecuteUnit_io_executeStage_inst_1_ex_tval_1),
    .io_executeStage_inst_1_ex_tval_2(ExecuteUnit_io_executeStage_inst_1_ex_tval_2),
    .io_executeStage_inst_1_ex_tval_12(ExecuteUnit_io_executeStage_inst_1_ex_tval_12),
    .io_executeStage_jump_branch_info_jump_regiser(ExecuteUnit_io_executeStage_jump_branch_info_jump_regiser),
    .io_executeStage_jump_branch_info_branch_inst(ExecuteUnit_io_executeStage_jump_branch_info_branch_inst),
    .io_executeStage_jump_branch_info_pred_branch(ExecuteUnit_io_executeStage_jump_branch_info_pred_branch),
    .io_executeStage_jump_branch_info_branch_target(ExecuteUnit_io_executeStage_jump_branch_info_branch_target),
    .io_executeStage_jump_branch_info_update_pht_index(ExecuteUnit_io_executeStage_jump_branch_info_update_pht_index),
    .io_csr_in_valid(ExecuteUnit_io_csr_in_valid),
    .io_csr_in_pc(ExecuteUnit_io_csr_in_pc),
    .io_csr_in_info_op(ExecuteUnit_io_csr_in_info_op),
    .io_csr_in_info_inst(ExecuteUnit_io_csr_in_info_inst),
    .io_csr_in_src_info_src1_data(ExecuteUnit_io_csr_in_src_info_src1_data),
    .io_csr_in_ex_exception_1(ExecuteUnit_io_csr_in_ex_exception_1),
    .io_csr_in_ex_exception_2(ExecuteUnit_io_csr_in_ex_exception_2),
    .io_csr_in_ex_exception_3(ExecuteUnit_io_csr_in_ex_exception_3),
    .io_csr_in_ex_exception_8(ExecuteUnit_io_csr_in_ex_exception_8),
    .io_csr_in_ex_exception_9(ExecuteUnit_io_csr_in_ex_exception_9),
    .io_csr_in_ex_exception_11(ExecuteUnit_io_csr_in_ex_exception_11),
    .io_csr_in_ex_exception_12(ExecuteUnit_io_csr_in_ex_exception_12),
    .io_csr_in_ex_interrupt_0(ExecuteUnit_io_csr_in_ex_interrupt_0),
    .io_csr_in_ex_interrupt_1(ExecuteUnit_io_csr_in_ex_interrupt_1),
    .io_csr_in_ex_interrupt_2(ExecuteUnit_io_csr_in_ex_interrupt_2),
    .io_csr_in_ex_interrupt_3(ExecuteUnit_io_csr_in_ex_interrupt_3),
    .io_csr_in_ex_interrupt_4(ExecuteUnit_io_csr_in_ex_interrupt_4),
    .io_csr_in_ex_interrupt_5(ExecuteUnit_io_csr_in_ex_interrupt_5),
    .io_csr_in_ex_interrupt_6(ExecuteUnit_io_csr_in_ex_interrupt_6),
    .io_csr_in_ex_interrupt_7(ExecuteUnit_io_csr_in_ex_interrupt_7),
    .io_csr_in_ex_interrupt_8(ExecuteUnit_io_csr_in_ex_interrupt_8),
    .io_csr_in_ex_interrupt_9(ExecuteUnit_io_csr_in_ex_interrupt_9),
    .io_csr_in_ex_interrupt_10(ExecuteUnit_io_csr_in_ex_interrupt_10),
    .io_csr_in_ex_interrupt_11(ExecuteUnit_io_csr_in_ex_interrupt_11),
    .io_csr_in_ex_tval_1(ExecuteUnit_io_csr_in_ex_tval_1),
    .io_csr_in_ex_tval_12(ExecuteUnit_io_csr_in_ex_tval_12),
    .io_csr_out_rdata(ExecuteUnit_io_csr_out_rdata),
    .io_csr_out_ex_exception_1(ExecuteUnit_io_csr_out_ex_exception_1),
    .io_csr_out_ex_exception_2(ExecuteUnit_io_csr_out_ex_exception_2),
    .io_csr_out_ex_exception_3(ExecuteUnit_io_csr_out_ex_exception_3),
    .io_csr_out_ex_exception_8(ExecuteUnit_io_csr_out_ex_exception_8),
    .io_csr_out_ex_exception_9(ExecuteUnit_io_csr_out_ex_exception_9),
    .io_csr_out_ex_exception_11(ExecuteUnit_io_csr_out_ex_exception_11),
    .io_csr_out_ex_exception_12(ExecuteUnit_io_csr_out_ex_exception_12),
    .io_csr_out_ex_interrupt_0(ExecuteUnit_io_csr_out_ex_interrupt_0),
    .io_csr_out_ex_interrupt_1(ExecuteUnit_io_csr_out_ex_interrupt_1),
    .io_csr_out_ex_interrupt_2(ExecuteUnit_io_csr_out_ex_interrupt_2),
    .io_csr_out_ex_interrupt_3(ExecuteUnit_io_csr_out_ex_interrupt_3),
    .io_csr_out_ex_interrupt_4(ExecuteUnit_io_csr_out_ex_interrupt_4),
    .io_csr_out_ex_interrupt_5(ExecuteUnit_io_csr_out_ex_interrupt_5),
    .io_csr_out_ex_interrupt_6(ExecuteUnit_io_csr_out_ex_interrupt_6),
    .io_csr_out_ex_interrupt_7(ExecuteUnit_io_csr_out_ex_interrupt_7),
    .io_csr_out_ex_interrupt_8(ExecuteUnit_io_csr_out_ex_interrupt_8),
    .io_csr_out_ex_interrupt_9(ExecuteUnit_io_csr_out_ex_interrupt_9),
    .io_csr_out_ex_interrupt_10(ExecuteUnit_io_csr_out_ex_interrupt_10),
    .io_csr_out_ex_interrupt_11(ExecuteUnit_io_csr_out_ex_interrupt_11),
    .io_csr_out_ex_tval_1(ExecuteUnit_io_csr_out_ex_tval_1),
    .io_csr_out_ex_tval_2(ExecuteUnit_io_csr_out_ex_tval_2),
    .io_csr_out_ex_tval_12(ExecuteUnit_io_csr_out_ex_tval_12),
    .io_csr_out_flush(ExecuteUnit_io_csr_out_flush),
    .io_csr_out_target(ExecuteUnit_io_csr_out_target),
    .io_bpu_pc(ExecuteUnit_io_bpu_pc),
    .io_bpu_update_pht_index(ExecuteUnit_io_bpu_update_pht_index),
    .io_bpu_branch_inst(ExecuteUnit_io_bpu_branch_inst),
    .io_bpu_branch(ExecuteUnit_io_bpu_branch),
    .io_fetchUnit_flush(ExecuteUnit_io_fetchUnit_flush),
    .io_fetchUnit_target(ExecuteUnit_io_fetchUnit_target),
    .io_decodeUnit_forward_0_exe_wen(ExecuteUnit_io_decodeUnit_forward_0_exe_wen),
    .io_decodeUnit_forward_0_exe_waddr(ExecuteUnit_io_decodeUnit_forward_0_exe_waddr),
    .io_decodeUnit_forward_0_exe_wdata(ExecuteUnit_io_decodeUnit_forward_0_exe_wdata),
    .io_decodeUnit_forward_0_is_load(ExecuteUnit_io_decodeUnit_forward_0_is_load),
    .io_decodeUnit_forward_1_exe_wen(ExecuteUnit_io_decodeUnit_forward_1_exe_wen),
    .io_decodeUnit_forward_1_exe_waddr(ExecuteUnit_io_decodeUnit_forward_1_exe_waddr),
    .io_decodeUnit_forward_1_exe_wdata(ExecuteUnit_io_decodeUnit_forward_1_exe_wdata),
    .io_decodeUnit_forward_1_is_load(ExecuteUnit_io_decodeUnit_forward_1_is_load),
    .io_memoryStage_inst_0_pc(ExecuteUnit_io_memoryStage_inst_0_pc),
    .io_memoryStage_inst_0_info_valid(ExecuteUnit_io_memoryStage_inst_0_info_valid),
    .io_memoryStage_inst_0_info_fusel(ExecuteUnit_io_memoryStage_inst_0_info_fusel),
    .io_memoryStage_inst_0_info_op(ExecuteUnit_io_memoryStage_inst_0_info_op),
    .io_memoryStage_inst_0_info_reg_wen(ExecuteUnit_io_memoryStage_inst_0_info_reg_wen),
    .io_memoryStage_inst_0_info_reg_waddr(ExecuteUnit_io_memoryStage_inst_0_info_reg_waddr),
    .io_memoryStage_inst_0_info_imm(ExecuteUnit_io_memoryStage_inst_0_info_imm),
    .io_memoryStage_inst_0_info_inst(ExecuteUnit_io_memoryStage_inst_0_info_inst),
    .io_memoryStage_inst_0_rd_info_wdata_0(ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_0),
    .io_memoryStage_inst_0_rd_info_wdata_1(ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_1),
    .io_memoryStage_inst_0_rd_info_wdata_2(ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_2),
    .io_memoryStage_inst_0_rd_info_wdata_3(ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_3),
    .io_memoryStage_inst_0_rd_info_wdata_4(ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_4),
    .io_memoryStage_inst_0_rd_info_wdata_5(ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_5),
    .io_memoryStage_inst_0_src_info_src1_data(ExecuteUnit_io_memoryStage_inst_0_src_info_src1_data),
    .io_memoryStage_inst_0_src_info_src2_data(ExecuteUnit_io_memoryStage_inst_0_src_info_src2_data),
    .io_memoryStage_inst_0_ex_exception_0(ExecuteUnit_io_memoryStage_inst_0_ex_exception_0),
    .io_memoryStage_inst_0_ex_exception_1(ExecuteUnit_io_memoryStage_inst_0_ex_exception_1),
    .io_memoryStage_inst_0_ex_exception_2(ExecuteUnit_io_memoryStage_inst_0_ex_exception_2),
    .io_memoryStage_inst_0_ex_exception_3(ExecuteUnit_io_memoryStage_inst_0_ex_exception_3),
    .io_memoryStage_inst_0_ex_exception_8(ExecuteUnit_io_memoryStage_inst_0_ex_exception_8),
    .io_memoryStage_inst_0_ex_exception_9(ExecuteUnit_io_memoryStage_inst_0_ex_exception_9),
    .io_memoryStage_inst_0_ex_exception_11(ExecuteUnit_io_memoryStage_inst_0_ex_exception_11),
    .io_memoryStage_inst_0_ex_exception_12(ExecuteUnit_io_memoryStage_inst_0_ex_exception_12),
    .io_memoryStage_inst_0_ex_interrupt_0(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_0),
    .io_memoryStage_inst_0_ex_interrupt_1(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_1),
    .io_memoryStage_inst_0_ex_interrupt_2(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_2),
    .io_memoryStage_inst_0_ex_interrupt_3(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_3),
    .io_memoryStage_inst_0_ex_interrupt_4(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_4),
    .io_memoryStage_inst_0_ex_interrupt_5(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_5),
    .io_memoryStage_inst_0_ex_interrupt_6(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_6),
    .io_memoryStage_inst_0_ex_interrupt_7(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_7),
    .io_memoryStage_inst_0_ex_interrupt_8(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_8),
    .io_memoryStage_inst_0_ex_interrupt_9(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_9),
    .io_memoryStage_inst_0_ex_interrupt_10(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_10),
    .io_memoryStage_inst_0_ex_interrupt_11(ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_11),
    .io_memoryStage_inst_0_ex_tval_0(ExecuteUnit_io_memoryStage_inst_0_ex_tval_0),
    .io_memoryStage_inst_0_ex_tval_1(ExecuteUnit_io_memoryStage_inst_0_ex_tval_1),
    .io_memoryStage_inst_0_ex_tval_2(ExecuteUnit_io_memoryStage_inst_0_ex_tval_2),
    .io_memoryStage_inst_0_ex_tval_12(ExecuteUnit_io_memoryStage_inst_0_ex_tval_12),
    .io_memoryStage_inst_1_pc(ExecuteUnit_io_memoryStage_inst_1_pc),
    .io_memoryStage_inst_1_info_valid(ExecuteUnit_io_memoryStage_inst_1_info_valid),
    .io_memoryStage_inst_1_info_fusel(ExecuteUnit_io_memoryStage_inst_1_info_fusel),
    .io_memoryStage_inst_1_info_op(ExecuteUnit_io_memoryStage_inst_1_info_op),
    .io_memoryStage_inst_1_info_reg_wen(ExecuteUnit_io_memoryStage_inst_1_info_reg_wen),
    .io_memoryStage_inst_1_info_reg_waddr(ExecuteUnit_io_memoryStage_inst_1_info_reg_waddr),
    .io_memoryStage_inst_1_info_imm(ExecuteUnit_io_memoryStage_inst_1_info_imm),
    .io_memoryStage_inst_1_info_inst(ExecuteUnit_io_memoryStage_inst_1_info_inst),
    .io_memoryStage_inst_1_rd_info_wdata_0(ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_0),
    .io_memoryStage_inst_1_rd_info_wdata_1(ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_1),
    .io_memoryStage_inst_1_rd_info_wdata_2(ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_2),
    .io_memoryStage_inst_1_rd_info_wdata_3(ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_3),
    .io_memoryStage_inst_1_rd_info_wdata_4(ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_4),
    .io_memoryStage_inst_1_rd_info_wdata_5(ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_5),
    .io_memoryStage_inst_1_src_info_src1_data(ExecuteUnit_io_memoryStage_inst_1_src_info_src1_data),
    .io_memoryStage_inst_1_src_info_src2_data(ExecuteUnit_io_memoryStage_inst_1_src_info_src2_data),
    .io_memoryStage_inst_1_ex_exception_0(ExecuteUnit_io_memoryStage_inst_1_ex_exception_0),
    .io_memoryStage_inst_1_ex_exception_1(ExecuteUnit_io_memoryStage_inst_1_ex_exception_1),
    .io_memoryStage_inst_1_ex_exception_2(ExecuteUnit_io_memoryStage_inst_1_ex_exception_2),
    .io_memoryStage_inst_1_ex_exception_3(ExecuteUnit_io_memoryStage_inst_1_ex_exception_3),
    .io_memoryStage_inst_1_ex_exception_8(ExecuteUnit_io_memoryStage_inst_1_ex_exception_8),
    .io_memoryStage_inst_1_ex_exception_9(ExecuteUnit_io_memoryStage_inst_1_ex_exception_9),
    .io_memoryStage_inst_1_ex_exception_11(ExecuteUnit_io_memoryStage_inst_1_ex_exception_11),
    .io_memoryStage_inst_1_ex_exception_12(ExecuteUnit_io_memoryStage_inst_1_ex_exception_12),
    .io_memoryStage_inst_1_ex_interrupt_0(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_0),
    .io_memoryStage_inst_1_ex_interrupt_1(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_1),
    .io_memoryStage_inst_1_ex_interrupt_2(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_2),
    .io_memoryStage_inst_1_ex_interrupt_3(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_3),
    .io_memoryStage_inst_1_ex_interrupt_4(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_4),
    .io_memoryStage_inst_1_ex_interrupt_5(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_5),
    .io_memoryStage_inst_1_ex_interrupt_6(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_6),
    .io_memoryStage_inst_1_ex_interrupt_7(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_7),
    .io_memoryStage_inst_1_ex_interrupt_8(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_8),
    .io_memoryStage_inst_1_ex_interrupt_9(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_9),
    .io_memoryStage_inst_1_ex_interrupt_10(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_10),
    .io_memoryStage_inst_1_ex_interrupt_11(ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_11),
    .io_memoryStage_inst_1_ex_tval_0(ExecuteUnit_io_memoryStage_inst_1_ex_tval_0),
    .io_memoryStage_inst_1_ex_tval_1(ExecuteUnit_io_memoryStage_inst_1_ex_tval_1),
    .io_memoryStage_inst_1_ex_tval_2(ExecuteUnit_io_memoryStage_inst_1_ex_tval_2),
    .io_memoryStage_inst_1_ex_tval_12(ExecuteUnit_io_memoryStage_inst_1_ex_tval_12),
    .io_dataMemory_addr(ExecuteUnit_io_dataMemory_addr)
  );
  Csr Csr ( // @[playground/src/Core.scala 33:30]
    .clock(Csr_clock),
    .reset(Csr_reset),
    .io_ext_int_ei(Csr_io_ext_int_ei),
    .io_ext_int_ti(Csr_io_ext_int_ti),
    .io_ext_int_si(Csr_io_ext_int_si),
    .io_decodeUnit_mode(Csr_io_decodeUnit_mode),
    .io_decodeUnit_interrupt(Csr_io_decodeUnit_interrupt),
    .io_executeUnit_in_valid(Csr_io_executeUnit_in_valid),
    .io_executeUnit_in_pc(Csr_io_executeUnit_in_pc),
    .io_executeUnit_in_info_op(Csr_io_executeUnit_in_info_op),
    .io_executeUnit_in_info_inst(Csr_io_executeUnit_in_info_inst),
    .io_executeUnit_in_src_info_src1_data(Csr_io_executeUnit_in_src_info_src1_data),
    .io_executeUnit_in_ex_exception_1(Csr_io_executeUnit_in_ex_exception_1),
    .io_executeUnit_in_ex_exception_2(Csr_io_executeUnit_in_ex_exception_2),
    .io_executeUnit_in_ex_exception_3(Csr_io_executeUnit_in_ex_exception_3),
    .io_executeUnit_in_ex_exception_8(Csr_io_executeUnit_in_ex_exception_8),
    .io_executeUnit_in_ex_exception_9(Csr_io_executeUnit_in_ex_exception_9),
    .io_executeUnit_in_ex_exception_11(Csr_io_executeUnit_in_ex_exception_11),
    .io_executeUnit_in_ex_exception_12(Csr_io_executeUnit_in_ex_exception_12),
    .io_executeUnit_in_ex_interrupt_0(Csr_io_executeUnit_in_ex_interrupt_0),
    .io_executeUnit_in_ex_interrupt_1(Csr_io_executeUnit_in_ex_interrupt_1),
    .io_executeUnit_in_ex_interrupt_2(Csr_io_executeUnit_in_ex_interrupt_2),
    .io_executeUnit_in_ex_interrupt_3(Csr_io_executeUnit_in_ex_interrupt_3),
    .io_executeUnit_in_ex_interrupt_4(Csr_io_executeUnit_in_ex_interrupt_4),
    .io_executeUnit_in_ex_interrupt_5(Csr_io_executeUnit_in_ex_interrupt_5),
    .io_executeUnit_in_ex_interrupt_6(Csr_io_executeUnit_in_ex_interrupt_6),
    .io_executeUnit_in_ex_interrupt_7(Csr_io_executeUnit_in_ex_interrupt_7),
    .io_executeUnit_in_ex_interrupt_8(Csr_io_executeUnit_in_ex_interrupt_8),
    .io_executeUnit_in_ex_interrupt_9(Csr_io_executeUnit_in_ex_interrupt_9),
    .io_executeUnit_in_ex_interrupt_10(Csr_io_executeUnit_in_ex_interrupt_10),
    .io_executeUnit_in_ex_interrupt_11(Csr_io_executeUnit_in_ex_interrupt_11),
    .io_executeUnit_in_ex_tval_1(Csr_io_executeUnit_in_ex_tval_1),
    .io_executeUnit_in_ex_tval_12(Csr_io_executeUnit_in_ex_tval_12),
    .io_executeUnit_out_rdata(Csr_io_executeUnit_out_rdata),
    .io_executeUnit_out_ex_exception_1(Csr_io_executeUnit_out_ex_exception_1),
    .io_executeUnit_out_ex_exception_2(Csr_io_executeUnit_out_ex_exception_2),
    .io_executeUnit_out_ex_exception_3(Csr_io_executeUnit_out_ex_exception_3),
    .io_executeUnit_out_ex_exception_8(Csr_io_executeUnit_out_ex_exception_8),
    .io_executeUnit_out_ex_exception_9(Csr_io_executeUnit_out_ex_exception_9),
    .io_executeUnit_out_ex_exception_11(Csr_io_executeUnit_out_ex_exception_11),
    .io_executeUnit_out_ex_exception_12(Csr_io_executeUnit_out_ex_exception_12),
    .io_executeUnit_out_ex_interrupt_0(Csr_io_executeUnit_out_ex_interrupt_0),
    .io_executeUnit_out_ex_interrupt_1(Csr_io_executeUnit_out_ex_interrupt_1),
    .io_executeUnit_out_ex_interrupt_2(Csr_io_executeUnit_out_ex_interrupt_2),
    .io_executeUnit_out_ex_interrupt_3(Csr_io_executeUnit_out_ex_interrupt_3),
    .io_executeUnit_out_ex_interrupt_4(Csr_io_executeUnit_out_ex_interrupt_4),
    .io_executeUnit_out_ex_interrupt_5(Csr_io_executeUnit_out_ex_interrupt_5),
    .io_executeUnit_out_ex_interrupt_6(Csr_io_executeUnit_out_ex_interrupt_6),
    .io_executeUnit_out_ex_interrupt_7(Csr_io_executeUnit_out_ex_interrupt_7),
    .io_executeUnit_out_ex_interrupt_8(Csr_io_executeUnit_out_ex_interrupt_8),
    .io_executeUnit_out_ex_interrupt_9(Csr_io_executeUnit_out_ex_interrupt_9),
    .io_executeUnit_out_ex_interrupt_10(Csr_io_executeUnit_out_ex_interrupt_10),
    .io_executeUnit_out_ex_interrupt_11(Csr_io_executeUnit_out_ex_interrupt_11),
    .io_executeUnit_out_ex_tval_1(Csr_io_executeUnit_out_ex_tval_1),
    .io_executeUnit_out_ex_tval_2(Csr_io_executeUnit_out_ex_tval_2),
    .io_executeUnit_out_ex_tval_12(Csr_io_executeUnit_out_ex_tval_12),
    .io_executeUnit_out_flush(Csr_io_executeUnit_out_flush),
    .io_executeUnit_out_target(Csr_io_executeUnit_out_target),
    .io_memoryUnit_in_pc(Csr_io_memoryUnit_in_pc),
    .io_memoryUnit_in_ex_exception_0(Csr_io_memoryUnit_in_ex_exception_0),
    .io_memoryUnit_in_ex_exception_1(Csr_io_memoryUnit_in_ex_exception_1),
    .io_memoryUnit_in_ex_exception_2(Csr_io_memoryUnit_in_ex_exception_2),
    .io_memoryUnit_in_ex_exception_3(Csr_io_memoryUnit_in_ex_exception_3),
    .io_memoryUnit_in_ex_exception_4(Csr_io_memoryUnit_in_ex_exception_4),
    .io_memoryUnit_in_ex_exception_5(Csr_io_memoryUnit_in_ex_exception_5),
    .io_memoryUnit_in_ex_exception_6(Csr_io_memoryUnit_in_ex_exception_6),
    .io_memoryUnit_in_ex_exception_7(Csr_io_memoryUnit_in_ex_exception_7),
    .io_memoryUnit_in_ex_exception_8(Csr_io_memoryUnit_in_ex_exception_8),
    .io_memoryUnit_in_ex_exception_9(Csr_io_memoryUnit_in_ex_exception_9),
    .io_memoryUnit_in_ex_exception_10(Csr_io_memoryUnit_in_ex_exception_10),
    .io_memoryUnit_in_ex_exception_11(Csr_io_memoryUnit_in_ex_exception_11),
    .io_memoryUnit_in_ex_exception_12(Csr_io_memoryUnit_in_ex_exception_12),
    .io_memoryUnit_in_ex_exception_13(Csr_io_memoryUnit_in_ex_exception_13),
    .io_memoryUnit_in_ex_exception_14(Csr_io_memoryUnit_in_ex_exception_14),
    .io_memoryUnit_in_ex_exception_15(Csr_io_memoryUnit_in_ex_exception_15),
    .io_memoryUnit_in_ex_interrupt_0(Csr_io_memoryUnit_in_ex_interrupt_0),
    .io_memoryUnit_in_ex_interrupt_1(Csr_io_memoryUnit_in_ex_interrupt_1),
    .io_memoryUnit_in_ex_interrupt_2(Csr_io_memoryUnit_in_ex_interrupt_2),
    .io_memoryUnit_in_ex_interrupt_3(Csr_io_memoryUnit_in_ex_interrupt_3),
    .io_memoryUnit_in_ex_interrupt_4(Csr_io_memoryUnit_in_ex_interrupt_4),
    .io_memoryUnit_in_ex_interrupt_5(Csr_io_memoryUnit_in_ex_interrupt_5),
    .io_memoryUnit_in_ex_interrupt_6(Csr_io_memoryUnit_in_ex_interrupt_6),
    .io_memoryUnit_in_ex_interrupt_7(Csr_io_memoryUnit_in_ex_interrupt_7),
    .io_memoryUnit_in_ex_interrupt_8(Csr_io_memoryUnit_in_ex_interrupt_8),
    .io_memoryUnit_in_ex_interrupt_9(Csr_io_memoryUnit_in_ex_interrupt_9),
    .io_memoryUnit_in_ex_interrupt_10(Csr_io_memoryUnit_in_ex_interrupt_10),
    .io_memoryUnit_in_ex_interrupt_11(Csr_io_memoryUnit_in_ex_interrupt_11),
    .io_memoryUnit_in_ex_tval_0(Csr_io_memoryUnit_in_ex_tval_0),
    .io_memoryUnit_in_ex_tval_1(Csr_io_memoryUnit_in_ex_tval_1),
    .io_memoryUnit_in_ex_tval_2(Csr_io_memoryUnit_in_ex_tval_2),
    .io_memoryUnit_in_ex_tval_3(Csr_io_memoryUnit_in_ex_tval_3),
    .io_memoryUnit_in_ex_tval_4(Csr_io_memoryUnit_in_ex_tval_4),
    .io_memoryUnit_in_ex_tval_5(Csr_io_memoryUnit_in_ex_tval_5),
    .io_memoryUnit_in_ex_tval_6(Csr_io_memoryUnit_in_ex_tval_6),
    .io_memoryUnit_in_ex_tval_7(Csr_io_memoryUnit_in_ex_tval_7),
    .io_memoryUnit_in_ex_tval_8(Csr_io_memoryUnit_in_ex_tval_8),
    .io_memoryUnit_in_ex_tval_9(Csr_io_memoryUnit_in_ex_tval_9),
    .io_memoryUnit_in_ex_tval_10(Csr_io_memoryUnit_in_ex_tval_10),
    .io_memoryUnit_in_ex_tval_11(Csr_io_memoryUnit_in_ex_tval_11),
    .io_memoryUnit_in_ex_tval_12(Csr_io_memoryUnit_in_ex_tval_12),
    .io_memoryUnit_in_ex_tval_13(Csr_io_memoryUnit_in_ex_tval_13),
    .io_memoryUnit_in_ex_tval_14(Csr_io_memoryUnit_in_ex_tval_14),
    .io_memoryUnit_in_ex_tval_15(Csr_io_memoryUnit_in_ex_tval_15),
    .io_memoryUnit_in_info_valid(Csr_io_memoryUnit_in_info_valid),
    .io_memoryUnit_in_info_fusel(Csr_io_memoryUnit_in_info_fusel),
    .io_memoryUnit_in_info_op(Csr_io_memoryUnit_in_info_op),
    .io_memoryUnit_in_lr_wen(Csr_io_memoryUnit_in_lr_wen),
    .io_memoryUnit_in_lr_wbit(Csr_io_memoryUnit_in_lr_wbit),
    .io_memoryUnit_in_lr_waddr(Csr_io_memoryUnit_in_lr_waddr),
    .io_memoryUnit_out_flush(Csr_io_memoryUnit_out_flush),
    .io_memoryUnit_out_target(Csr_io_memoryUnit_out_target),
    .io_memoryUnit_out_lr(Csr_io_memoryUnit_out_lr),
    .io_memoryUnit_out_lr_addr(Csr_io_memoryUnit_out_lr_addr),
    .io_tlb_satp(Csr_io_tlb_satp),
    .io_tlb_mstatus(Csr_io_tlb_mstatus),
    .io_tlb_imode(Csr_io_tlb_imode),
    .io_tlb_dmode(Csr_io_tlb_dmode)
  );
  MemoryStage MemoryStage ( // @[playground/src/Core.scala 34:30]
    .clock(MemoryStage_clock),
    .reset(MemoryStage_reset),
    .io_ctrl_allow_to_go(MemoryStage_io_ctrl_allow_to_go),
    .io_ctrl_clear(MemoryStage_io_ctrl_clear),
    .io_executeUnit_inst_0_pc(MemoryStage_io_executeUnit_inst_0_pc),
    .io_executeUnit_inst_0_info_valid(MemoryStage_io_executeUnit_inst_0_info_valid),
    .io_executeUnit_inst_0_info_fusel(MemoryStage_io_executeUnit_inst_0_info_fusel),
    .io_executeUnit_inst_0_info_op(MemoryStage_io_executeUnit_inst_0_info_op),
    .io_executeUnit_inst_0_info_reg_wen(MemoryStage_io_executeUnit_inst_0_info_reg_wen),
    .io_executeUnit_inst_0_info_reg_waddr(MemoryStage_io_executeUnit_inst_0_info_reg_waddr),
    .io_executeUnit_inst_0_info_imm(MemoryStage_io_executeUnit_inst_0_info_imm),
    .io_executeUnit_inst_0_info_inst(MemoryStage_io_executeUnit_inst_0_info_inst),
    .io_executeUnit_inst_0_rd_info_wdata_0(MemoryStage_io_executeUnit_inst_0_rd_info_wdata_0),
    .io_executeUnit_inst_0_rd_info_wdata_2(MemoryStage_io_executeUnit_inst_0_rd_info_wdata_2),
    .io_executeUnit_inst_0_rd_info_wdata_3(MemoryStage_io_executeUnit_inst_0_rd_info_wdata_3),
    .io_executeUnit_inst_0_rd_info_wdata_5(MemoryStage_io_executeUnit_inst_0_rd_info_wdata_5),
    .io_executeUnit_inst_0_src_info_src1_data(MemoryStage_io_executeUnit_inst_0_src_info_src1_data),
    .io_executeUnit_inst_0_src_info_src2_data(MemoryStage_io_executeUnit_inst_0_src_info_src2_data),
    .io_executeUnit_inst_0_ex_exception_0(MemoryStage_io_executeUnit_inst_0_ex_exception_0),
    .io_executeUnit_inst_0_ex_exception_1(MemoryStage_io_executeUnit_inst_0_ex_exception_1),
    .io_executeUnit_inst_0_ex_exception_2(MemoryStage_io_executeUnit_inst_0_ex_exception_2),
    .io_executeUnit_inst_0_ex_exception_3(MemoryStage_io_executeUnit_inst_0_ex_exception_3),
    .io_executeUnit_inst_0_ex_exception_8(MemoryStage_io_executeUnit_inst_0_ex_exception_8),
    .io_executeUnit_inst_0_ex_exception_9(MemoryStage_io_executeUnit_inst_0_ex_exception_9),
    .io_executeUnit_inst_0_ex_exception_11(MemoryStage_io_executeUnit_inst_0_ex_exception_11),
    .io_executeUnit_inst_0_ex_exception_12(MemoryStage_io_executeUnit_inst_0_ex_exception_12),
    .io_executeUnit_inst_0_ex_interrupt_0(MemoryStage_io_executeUnit_inst_0_ex_interrupt_0),
    .io_executeUnit_inst_0_ex_interrupt_1(MemoryStage_io_executeUnit_inst_0_ex_interrupt_1),
    .io_executeUnit_inst_0_ex_interrupt_2(MemoryStage_io_executeUnit_inst_0_ex_interrupt_2),
    .io_executeUnit_inst_0_ex_interrupt_3(MemoryStage_io_executeUnit_inst_0_ex_interrupt_3),
    .io_executeUnit_inst_0_ex_interrupt_4(MemoryStage_io_executeUnit_inst_0_ex_interrupt_4),
    .io_executeUnit_inst_0_ex_interrupt_5(MemoryStage_io_executeUnit_inst_0_ex_interrupt_5),
    .io_executeUnit_inst_0_ex_interrupt_6(MemoryStage_io_executeUnit_inst_0_ex_interrupt_6),
    .io_executeUnit_inst_0_ex_interrupt_7(MemoryStage_io_executeUnit_inst_0_ex_interrupt_7),
    .io_executeUnit_inst_0_ex_interrupt_8(MemoryStage_io_executeUnit_inst_0_ex_interrupt_8),
    .io_executeUnit_inst_0_ex_interrupt_9(MemoryStage_io_executeUnit_inst_0_ex_interrupt_9),
    .io_executeUnit_inst_0_ex_interrupt_10(MemoryStage_io_executeUnit_inst_0_ex_interrupt_10),
    .io_executeUnit_inst_0_ex_interrupt_11(MemoryStage_io_executeUnit_inst_0_ex_interrupt_11),
    .io_executeUnit_inst_0_ex_tval_0(MemoryStage_io_executeUnit_inst_0_ex_tval_0),
    .io_executeUnit_inst_0_ex_tval_1(MemoryStage_io_executeUnit_inst_0_ex_tval_1),
    .io_executeUnit_inst_0_ex_tval_2(MemoryStage_io_executeUnit_inst_0_ex_tval_2),
    .io_executeUnit_inst_0_ex_tval_12(MemoryStage_io_executeUnit_inst_0_ex_tval_12),
    .io_executeUnit_inst_1_pc(MemoryStage_io_executeUnit_inst_1_pc),
    .io_executeUnit_inst_1_info_valid(MemoryStage_io_executeUnit_inst_1_info_valid),
    .io_executeUnit_inst_1_info_fusel(MemoryStage_io_executeUnit_inst_1_info_fusel),
    .io_executeUnit_inst_1_info_op(MemoryStage_io_executeUnit_inst_1_info_op),
    .io_executeUnit_inst_1_info_reg_wen(MemoryStage_io_executeUnit_inst_1_info_reg_wen),
    .io_executeUnit_inst_1_info_reg_waddr(MemoryStage_io_executeUnit_inst_1_info_reg_waddr),
    .io_executeUnit_inst_1_info_imm(MemoryStage_io_executeUnit_inst_1_info_imm),
    .io_executeUnit_inst_1_info_inst(MemoryStage_io_executeUnit_inst_1_info_inst),
    .io_executeUnit_inst_1_rd_info_wdata_0(MemoryStage_io_executeUnit_inst_1_rd_info_wdata_0),
    .io_executeUnit_inst_1_rd_info_wdata_2(MemoryStage_io_executeUnit_inst_1_rd_info_wdata_2),
    .io_executeUnit_inst_1_rd_info_wdata_3(MemoryStage_io_executeUnit_inst_1_rd_info_wdata_3),
    .io_executeUnit_inst_1_rd_info_wdata_5(MemoryStage_io_executeUnit_inst_1_rd_info_wdata_5),
    .io_executeUnit_inst_1_src_info_src1_data(MemoryStage_io_executeUnit_inst_1_src_info_src1_data),
    .io_executeUnit_inst_1_src_info_src2_data(MemoryStage_io_executeUnit_inst_1_src_info_src2_data),
    .io_executeUnit_inst_1_ex_exception_0(MemoryStage_io_executeUnit_inst_1_ex_exception_0),
    .io_executeUnit_inst_1_ex_exception_1(MemoryStage_io_executeUnit_inst_1_ex_exception_1),
    .io_executeUnit_inst_1_ex_exception_2(MemoryStage_io_executeUnit_inst_1_ex_exception_2),
    .io_executeUnit_inst_1_ex_exception_3(MemoryStage_io_executeUnit_inst_1_ex_exception_3),
    .io_executeUnit_inst_1_ex_exception_8(MemoryStage_io_executeUnit_inst_1_ex_exception_8),
    .io_executeUnit_inst_1_ex_exception_9(MemoryStage_io_executeUnit_inst_1_ex_exception_9),
    .io_executeUnit_inst_1_ex_exception_11(MemoryStage_io_executeUnit_inst_1_ex_exception_11),
    .io_executeUnit_inst_1_ex_exception_12(MemoryStage_io_executeUnit_inst_1_ex_exception_12),
    .io_executeUnit_inst_1_ex_interrupt_0(MemoryStage_io_executeUnit_inst_1_ex_interrupt_0),
    .io_executeUnit_inst_1_ex_interrupt_1(MemoryStage_io_executeUnit_inst_1_ex_interrupt_1),
    .io_executeUnit_inst_1_ex_interrupt_2(MemoryStage_io_executeUnit_inst_1_ex_interrupt_2),
    .io_executeUnit_inst_1_ex_interrupt_3(MemoryStage_io_executeUnit_inst_1_ex_interrupt_3),
    .io_executeUnit_inst_1_ex_interrupt_4(MemoryStage_io_executeUnit_inst_1_ex_interrupt_4),
    .io_executeUnit_inst_1_ex_interrupt_5(MemoryStage_io_executeUnit_inst_1_ex_interrupt_5),
    .io_executeUnit_inst_1_ex_interrupt_6(MemoryStage_io_executeUnit_inst_1_ex_interrupt_6),
    .io_executeUnit_inst_1_ex_interrupt_7(MemoryStage_io_executeUnit_inst_1_ex_interrupt_7),
    .io_executeUnit_inst_1_ex_interrupt_8(MemoryStage_io_executeUnit_inst_1_ex_interrupt_8),
    .io_executeUnit_inst_1_ex_interrupt_9(MemoryStage_io_executeUnit_inst_1_ex_interrupt_9),
    .io_executeUnit_inst_1_ex_interrupt_10(MemoryStage_io_executeUnit_inst_1_ex_interrupt_10),
    .io_executeUnit_inst_1_ex_interrupt_11(MemoryStage_io_executeUnit_inst_1_ex_interrupt_11),
    .io_executeUnit_inst_1_ex_tval_0(MemoryStage_io_executeUnit_inst_1_ex_tval_0),
    .io_executeUnit_inst_1_ex_tval_1(MemoryStage_io_executeUnit_inst_1_ex_tval_1),
    .io_executeUnit_inst_1_ex_tval_2(MemoryStage_io_executeUnit_inst_1_ex_tval_2),
    .io_executeUnit_inst_1_ex_tval_12(MemoryStage_io_executeUnit_inst_1_ex_tval_12),
    .io_memoryUnit_inst_0_pc(MemoryStage_io_memoryUnit_inst_0_pc),
    .io_memoryUnit_inst_0_info_valid(MemoryStage_io_memoryUnit_inst_0_info_valid),
    .io_memoryUnit_inst_0_info_fusel(MemoryStage_io_memoryUnit_inst_0_info_fusel),
    .io_memoryUnit_inst_0_info_op(MemoryStage_io_memoryUnit_inst_0_info_op),
    .io_memoryUnit_inst_0_info_reg_wen(MemoryStage_io_memoryUnit_inst_0_info_reg_wen),
    .io_memoryUnit_inst_0_info_reg_waddr(MemoryStage_io_memoryUnit_inst_0_info_reg_waddr),
    .io_memoryUnit_inst_0_info_imm(MemoryStage_io_memoryUnit_inst_0_info_imm),
    .io_memoryUnit_inst_0_info_inst(MemoryStage_io_memoryUnit_inst_0_info_inst),
    .io_memoryUnit_inst_0_rd_info_wdata_0(MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_0),
    .io_memoryUnit_inst_0_rd_info_wdata_2(MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_2),
    .io_memoryUnit_inst_0_rd_info_wdata_3(MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_3),
    .io_memoryUnit_inst_0_rd_info_wdata_5(MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_5),
    .io_memoryUnit_inst_0_src_info_src1_data(MemoryStage_io_memoryUnit_inst_0_src_info_src1_data),
    .io_memoryUnit_inst_0_src_info_src2_data(MemoryStage_io_memoryUnit_inst_0_src_info_src2_data),
    .io_memoryUnit_inst_0_ex_exception_0(MemoryStage_io_memoryUnit_inst_0_ex_exception_0),
    .io_memoryUnit_inst_0_ex_exception_1(MemoryStage_io_memoryUnit_inst_0_ex_exception_1),
    .io_memoryUnit_inst_0_ex_exception_2(MemoryStage_io_memoryUnit_inst_0_ex_exception_2),
    .io_memoryUnit_inst_0_ex_exception_3(MemoryStage_io_memoryUnit_inst_0_ex_exception_3),
    .io_memoryUnit_inst_0_ex_exception_8(MemoryStage_io_memoryUnit_inst_0_ex_exception_8),
    .io_memoryUnit_inst_0_ex_exception_9(MemoryStage_io_memoryUnit_inst_0_ex_exception_9),
    .io_memoryUnit_inst_0_ex_exception_11(MemoryStage_io_memoryUnit_inst_0_ex_exception_11),
    .io_memoryUnit_inst_0_ex_exception_12(MemoryStage_io_memoryUnit_inst_0_ex_exception_12),
    .io_memoryUnit_inst_0_ex_interrupt_0(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_0),
    .io_memoryUnit_inst_0_ex_interrupt_1(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_1),
    .io_memoryUnit_inst_0_ex_interrupt_2(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_2),
    .io_memoryUnit_inst_0_ex_interrupt_3(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_3),
    .io_memoryUnit_inst_0_ex_interrupt_4(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_4),
    .io_memoryUnit_inst_0_ex_interrupt_5(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_5),
    .io_memoryUnit_inst_0_ex_interrupt_6(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_6),
    .io_memoryUnit_inst_0_ex_interrupt_7(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_7),
    .io_memoryUnit_inst_0_ex_interrupt_8(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_8),
    .io_memoryUnit_inst_0_ex_interrupt_9(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_9),
    .io_memoryUnit_inst_0_ex_interrupt_10(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_10),
    .io_memoryUnit_inst_0_ex_interrupt_11(MemoryStage_io_memoryUnit_inst_0_ex_interrupt_11),
    .io_memoryUnit_inst_0_ex_tval_0(MemoryStage_io_memoryUnit_inst_0_ex_tval_0),
    .io_memoryUnit_inst_0_ex_tval_1(MemoryStage_io_memoryUnit_inst_0_ex_tval_1),
    .io_memoryUnit_inst_0_ex_tval_2(MemoryStage_io_memoryUnit_inst_0_ex_tval_2),
    .io_memoryUnit_inst_0_ex_tval_12(MemoryStage_io_memoryUnit_inst_0_ex_tval_12),
    .io_memoryUnit_inst_1_pc(MemoryStage_io_memoryUnit_inst_1_pc),
    .io_memoryUnit_inst_1_info_valid(MemoryStage_io_memoryUnit_inst_1_info_valid),
    .io_memoryUnit_inst_1_info_fusel(MemoryStage_io_memoryUnit_inst_1_info_fusel),
    .io_memoryUnit_inst_1_info_op(MemoryStage_io_memoryUnit_inst_1_info_op),
    .io_memoryUnit_inst_1_info_reg_wen(MemoryStage_io_memoryUnit_inst_1_info_reg_wen),
    .io_memoryUnit_inst_1_info_reg_waddr(MemoryStage_io_memoryUnit_inst_1_info_reg_waddr),
    .io_memoryUnit_inst_1_info_imm(MemoryStage_io_memoryUnit_inst_1_info_imm),
    .io_memoryUnit_inst_1_info_inst(MemoryStage_io_memoryUnit_inst_1_info_inst),
    .io_memoryUnit_inst_1_rd_info_wdata_0(MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_0),
    .io_memoryUnit_inst_1_rd_info_wdata_2(MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_2),
    .io_memoryUnit_inst_1_rd_info_wdata_3(MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_3),
    .io_memoryUnit_inst_1_rd_info_wdata_5(MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_5),
    .io_memoryUnit_inst_1_src_info_src1_data(MemoryStage_io_memoryUnit_inst_1_src_info_src1_data),
    .io_memoryUnit_inst_1_src_info_src2_data(MemoryStage_io_memoryUnit_inst_1_src_info_src2_data),
    .io_memoryUnit_inst_1_ex_exception_0(MemoryStage_io_memoryUnit_inst_1_ex_exception_0),
    .io_memoryUnit_inst_1_ex_exception_1(MemoryStage_io_memoryUnit_inst_1_ex_exception_1),
    .io_memoryUnit_inst_1_ex_exception_2(MemoryStage_io_memoryUnit_inst_1_ex_exception_2),
    .io_memoryUnit_inst_1_ex_exception_3(MemoryStage_io_memoryUnit_inst_1_ex_exception_3),
    .io_memoryUnit_inst_1_ex_exception_8(MemoryStage_io_memoryUnit_inst_1_ex_exception_8),
    .io_memoryUnit_inst_1_ex_exception_9(MemoryStage_io_memoryUnit_inst_1_ex_exception_9),
    .io_memoryUnit_inst_1_ex_exception_11(MemoryStage_io_memoryUnit_inst_1_ex_exception_11),
    .io_memoryUnit_inst_1_ex_exception_12(MemoryStage_io_memoryUnit_inst_1_ex_exception_12),
    .io_memoryUnit_inst_1_ex_interrupt_0(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_0),
    .io_memoryUnit_inst_1_ex_interrupt_1(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_1),
    .io_memoryUnit_inst_1_ex_interrupt_2(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_2),
    .io_memoryUnit_inst_1_ex_interrupt_3(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_3),
    .io_memoryUnit_inst_1_ex_interrupt_4(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_4),
    .io_memoryUnit_inst_1_ex_interrupt_5(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_5),
    .io_memoryUnit_inst_1_ex_interrupt_6(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_6),
    .io_memoryUnit_inst_1_ex_interrupt_7(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_7),
    .io_memoryUnit_inst_1_ex_interrupt_8(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_8),
    .io_memoryUnit_inst_1_ex_interrupt_9(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_9),
    .io_memoryUnit_inst_1_ex_interrupt_10(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_10),
    .io_memoryUnit_inst_1_ex_interrupt_11(MemoryStage_io_memoryUnit_inst_1_ex_interrupt_11),
    .io_memoryUnit_inst_1_ex_tval_0(MemoryStage_io_memoryUnit_inst_1_ex_tval_0),
    .io_memoryUnit_inst_1_ex_tval_1(MemoryStage_io_memoryUnit_inst_1_ex_tval_1),
    .io_memoryUnit_inst_1_ex_tval_2(MemoryStage_io_memoryUnit_inst_1_ex_tval_2),
    .io_memoryUnit_inst_1_ex_tval_12(MemoryStage_io_memoryUnit_inst_1_ex_tval_12)
  );
  MemoryUnit MemoryUnit ( // @[playground/src/Core.scala 35:30]
    .clock(MemoryUnit_clock),
    .reset(MemoryUnit_reset),
    .io_ctrl_flush(MemoryUnit_io_ctrl_flush),
    .io_ctrl_mem_stall(MemoryUnit_io_ctrl_mem_stall),
    .io_ctrl_allow_to_go(MemoryUnit_io_ctrl_allow_to_go),
    .io_ctrl_fence_i(MemoryUnit_io_ctrl_fence_i),
    .io_ctrl_complete_single_request(MemoryUnit_io_ctrl_complete_single_request),
    .io_ctrl_sfence_vma_valid(MemoryUnit_io_ctrl_sfence_vma_valid),
    .io_ctrl_sfence_vma_src_info_src1_data(MemoryUnit_io_ctrl_sfence_vma_src_info_src1_data),
    .io_ctrl_sfence_vma_src_info_src2_data(MemoryUnit_io_ctrl_sfence_vma_src_info_src2_data),
    .io_memoryStage_inst_0_pc(MemoryUnit_io_memoryStage_inst_0_pc),
    .io_memoryStage_inst_0_info_valid(MemoryUnit_io_memoryStage_inst_0_info_valid),
    .io_memoryStage_inst_0_info_fusel(MemoryUnit_io_memoryStage_inst_0_info_fusel),
    .io_memoryStage_inst_0_info_op(MemoryUnit_io_memoryStage_inst_0_info_op),
    .io_memoryStage_inst_0_info_reg_wen(MemoryUnit_io_memoryStage_inst_0_info_reg_wen),
    .io_memoryStage_inst_0_info_reg_waddr(MemoryUnit_io_memoryStage_inst_0_info_reg_waddr),
    .io_memoryStage_inst_0_info_imm(MemoryUnit_io_memoryStage_inst_0_info_imm),
    .io_memoryStage_inst_0_info_inst(MemoryUnit_io_memoryStage_inst_0_info_inst),
    .io_memoryStage_inst_0_rd_info_wdata_0(MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_0),
    .io_memoryStage_inst_0_rd_info_wdata_2(MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_2),
    .io_memoryStage_inst_0_rd_info_wdata_3(MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_3),
    .io_memoryStage_inst_0_rd_info_wdata_5(MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_5),
    .io_memoryStage_inst_0_src_info_src1_data(MemoryUnit_io_memoryStage_inst_0_src_info_src1_data),
    .io_memoryStage_inst_0_src_info_src2_data(MemoryUnit_io_memoryStage_inst_0_src_info_src2_data),
    .io_memoryStage_inst_0_ex_exception_0(MemoryUnit_io_memoryStage_inst_0_ex_exception_0),
    .io_memoryStage_inst_0_ex_exception_1(MemoryUnit_io_memoryStage_inst_0_ex_exception_1),
    .io_memoryStage_inst_0_ex_exception_2(MemoryUnit_io_memoryStage_inst_0_ex_exception_2),
    .io_memoryStage_inst_0_ex_exception_3(MemoryUnit_io_memoryStage_inst_0_ex_exception_3),
    .io_memoryStage_inst_0_ex_exception_8(MemoryUnit_io_memoryStage_inst_0_ex_exception_8),
    .io_memoryStage_inst_0_ex_exception_9(MemoryUnit_io_memoryStage_inst_0_ex_exception_9),
    .io_memoryStage_inst_0_ex_exception_11(MemoryUnit_io_memoryStage_inst_0_ex_exception_11),
    .io_memoryStage_inst_0_ex_exception_12(MemoryUnit_io_memoryStage_inst_0_ex_exception_12),
    .io_memoryStage_inst_0_ex_interrupt_0(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_0),
    .io_memoryStage_inst_0_ex_interrupt_1(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_1),
    .io_memoryStage_inst_0_ex_interrupt_2(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_2),
    .io_memoryStage_inst_0_ex_interrupt_3(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_3),
    .io_memoryStage_inst_0_ex_interrupt_4(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_4),
    .io_memoryStage_inst_0_ex_interrupt_5(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_5),
    .io_memoryStage_inst_0_ex_interrupt_6(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_6),
    .io_memoryStage_inst_0_ex_interrupt_7(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_7),
    .io_memoryStage_inst_0_ex_interrupt_8(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_8),
    .io_memoryStage_inst_0_ex_interrupt_9(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_9),
    .io_memoryStage_inst_0_ex_interrupt_10(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_10),
    .io_memoryStage_inst_0_ex_interrupt_11(MemoryUnit_io_memoryStage_inst_0_ex_interrupt_11),
    .io_memoryStage_inst_0_ex_tval_0(MemoryUnit_io_memoryStage_inst_0_ex_tval_0),
    .io_memoryStage_inst_0_ex_tval_1(MemoryUnit_io_memoryStage_inst_0_ex_tval_1),
    .io_memoryStage_inst_0_ex_tval_2(MemoryUnit_io_memoryStage_inst_0_ex_tval_2),
    .io_memoryStage_inst_0_ex_tval_12(MemoryUnit_io_memoryStage_inst_0_ex_tval_12),
    .io_memoryStage_inst_1_pc(MemoryUnit_io_memoryStage_inst_1_pc),
    .io_memoryStage_inst_1_info_valid(MemoryUnit_io_memoryStage_inst_1_info_valid),
    .io_memoryStage_inst_1_info_fusel(MemoryUnit_io_memoryStage_inst_1_info_fusel),
    .io_memoryStage_inst_1_info_op(MemoryUnit_io_memoryStage_inst_1_info_op),
    .io_memoryStage_inst_1_info_reg_wen(MemoryUnit_io_memoryStage_inst_1_info_reg_wen),
    .io_memoryStage_inst_1_info_reg_waddr(MemoryUnit_io_memoryStage_inst_1_info_reg_waddr),
    .io_memoryStage_inst_1_info_imm(MemoryUnit_io_memoryStage_inst_1_info_imm),
    .io_memoryStage_inst_1_info_inst(MemoryUnit_io_memoryStage_inst_1_info_inst),
    .io_memoryStage_inst_1_rd_info_wdata_0(MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_0),
    .io_memoryStage_inst_1_rd_info_wdata_2(MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_2),
    .io_memoryStage_inst_1_rd_info_wdata_3(MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_3),
    .io_memoryStage_inst_1_rd_info_wdata_5(MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_5),
    .io_memoryStage_inst_1_src_info_src1_data(MemoryUnit_io_memoryStage_inst_1_src_info_src1_data),
    .io_memoryStage_inst_1_src_info_src2_data(MemoryUnit_io_memoryStage_inst_1_src_info_src2_data),
    .io_memoryStage_inst_1_ex_exception_0(MemoryUnit_io_memoryStage_inst_1_ex_exception_0),
    .io_memoryStage_inst_1_ex_exception_1(MemoryUnit_io_memoryStage_inst_1_ex_exception_1),
    .io_memoryStage_inst_1_ex_exception_2(MemoryUnit_io_memoryStage_inst_1_ex_exception_2),
    .io_memoryStage_inst_1_ex_exception_3(MemoryUnit_io_memoryStage_inst_1_ex_exception_3),
    .io_memoryStage_inst_1_ex_exception_8(MemoryUnit_io_memoryStage_inst_1_ex_exception_8),
    .io_memoryStage_inst_1_ex_exception_9(MemoryUnit_io_memoryStage_inst_1_ex_exception_9),
    .io_memoryStage_inst_1_ex_exception_11(MemoryUnit_io_memoryStage_inst_1_ex_exception_11),
    .io_memoryStage_inst_1_ex_exception_12(MemoryUnit_io_memoryStage_inst_1_ex_exception_12),
    .io_memoryStage_inst_1_ex_interrupt_0(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_0),
    .io_memoryStage_inst_1_ex_interrupt_1(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_1),
    .io_memoryStage_inst_1_ex_interrupt_2(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_2),
    .io_memoryStage_inst_1_ex_interrupt_3(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_3),
    .io_memoryStage_inst_1_ex_interrupt_4(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_4),
    .io_memoryStage_inst_1_ex_interrupt_5(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_5),
    .io_memoryStage_inst_1_ex_interrupt_6(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_6),
    .io_memoryStage_inst_1_ex_interrupt_7(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_7),
    .io_memoryStage_inst_1_ex_interrupt_8(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_8),
    .io_memoryStage_inst_1_ex_interrupt_9(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_9),
    .io_memoryStage_inst_1_ex_interrupt_10(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_10),
    .io_memoryStage_inst_1_ex_interrupt_11(MemoryUnit_io_memoryStage_inst_1_ex_interrupt_11),
    .io_memoryStage_inst_1_ex_tval_0(MemoryUnit_io_memoryStage_inst_1_ex_tval_0),
    .io_memoryStage_inst_1_ex_tval_1(MemoryUnit_io_memoryStage_inst_1_ex_tval_1),
    .io_memoryStage_inst_1_ex_tval_2(MemoryUnit_io_memoryStage_inst_1_ex_tval_2),
    .io_memoryStage_inst_1_ex_tval_12(MemoryUnit_io_memoryStage_inst_1_ex_tval_12),
    .io_fetchUnit_flush(MemoryUnit_io_fetchUnit_flush),
    .io_fetchUnit_target(MemoryUnit_io_fetchUnit_target),
    .io_decodeUnit_0_wen(MemoryUnit_io_decodeUnit_0_wen),
    .io_decodeUnit_0_waddr(MemoryUnit_io_decodeUnit_0_waddr),
    .io_decodeUnit_0_wdata(MemoryUnit_io_decodeUnit_0_wdata),
    .io_decodeUnit_1_wen(MemoryUnit_io_decodeUnit_1_wen),
    .io_decodeUnit_1_waddr(MemoryUnit_io_decodeUnit_1_waddr),
    .io_decodeUnit_1_wdata(MemoryUnit_io_decodeUnit_1_wdata),
    .io_csr_in_pc(MemoryUnit_io_csr_in_pc),
    .io_csr_in_ex_exception_0(MemoryUnit_io_csr_in_ex_exception_0),
    .io_csr_in_ex_exception_1(MemoryUnit_io_csr_in_ex_exception_1),
    .io_csr_in_ex_exception_2(MemoryUnit_io_csr_in_ex_exception_2),
    .io_csr_in_ex_exception_3(MemoryUnit_io_csr_in_ex_exception_3),
    .io_csr_in_ex_exception_4(MemoryUnit_io_csr_in_ex_exception_4),
    .io_csr_in_ex_exception_5(MemoryUnit_io_csr_in_ex_exception_5),
    .io_csr_in_ex_exception_6(MemoryUnit_io_csr_in_ex_exception_6),
    .io_csr_in_ex_exception_7(MemoryUnit_io_csr_in_ex_exception_7),
    .io_csr_in_ex_exception_8(MemoryUnit_io_csr_in_ex_exception_8),
    .io_csr_in_ex_exception_9(MemoryUnit_io_csr_in_ex_exception_9),
    .io_csr_in_ex_exception_10(MemoryUnit_io_csr_in_ex_exception_10),
    .io_csr_in_ex_exception_11(MemoryUnit_io_csr_in_ex_exception_11),
    .io_csr_in_ex_exception_12(MemoryUnit_io_csr_in_ex_exception_12),
    .io_csr_in_ex_exception_13(MemoryUnit_io_csr_in_ex_exception_13),
    .io_csr_in_ex_exception_14(MemoryUnit_io_csr_in_ex_exception_14),
    .io_csr_in_ex_exception_15(MemoryUnit_io_csr_in_ex_exception_15),
    .io_csr_in_ex_interrupt_0(MemoryUnit_io_csr_in_ex_interrupt_0),
    .io_csr_in_ex_interrupt_1(MemoryUnit_io_csr_in_ex_interrupt_1),
    .io_csr_in_ex_interrupt_2(MemoryUnit_io_csr_in_ex_interrupt_2),
    .io_csr_in_ex_interrupt_3(MemoryUnit_io_csr_in_ex_interrupt_3),
    .io_csr_in_ex_interrupt_4(MemoryUnit_io_csr_in_ex_interrupt_4),
    .io_csr_in_ex_interrupt_5(MemoryUnit_io_csr_in_ex_interrupt_5),
    .io_csr_in_ex_interrupt_6(MemoryUnit_io_csr_in_ex_interrupt_6),
    .io_csr_in_ex_interrupt_7(MemoryUnit_io_csr_in_ex_interrupt_7),
    .io_csr_in_ex_interrupt_8(MemoryUnit_io_csr_in_ex_interrupt_8),
    .io_csr_in_ex_interrupt_9(MemoryUnit_io_csr_in_ex_interrupt_9),
    .io_csr_in_ex_interrupt_10(MemoryUnit_io_csr_in_ex_interrupt_10),
    .io_csr_in_ex_interrupt_11(MemoryUnit_io_csr_in_ex_interrupt_11),
    .io_csr_in_ex_tval_0(MemoryUnit_io_csr_in_ex_tval_0),
    .io_csr_in_ex_tval_1(MemoryUnit_io_csr_in_ex_tval_1),
    .io_csr_in_ex_tval_2(MemoryUnit_io_csr_in_ex_tval_2),
    .io_csr_in_ex_tval_3(MemoryUnit_io_csr_in_ex_tval_3),
    .io_csr_in_ex_tval_4(MemoryUnit_io_csr_in_ex_tval_4),
    .io_csr_in_ex_tval_5(MemoryUnit_io_csr_in_ex_tval_5),
    .io_csr_in_ex_tval_6(MemoryUnit_io_csr_in_ex_tval_6),
    .io_csr_in_ex_tval_7(MemoryUnit_io_csr_in_ex_tval_7),
    .io_csr_in_ex_tval_8(MemoryUnit_io_csr_in_ex_tval_8),
    .io_csr_in_ex_tval_9(MemoryUnit_io_csr_in_ex_tval_9),
    .io_csr_in_ex_tval_10(MemoryUnit_io_csr_in_ex_tval_10),
    .io_csr_in_ex_tval_11(MemoryUnit_io_csr_in_ex_tval_11),
    .io_csr_in_ex_tval_12(MemoryUnit_io_csr_in_ex_tval_12),
    .io_csr_in_ex_tval_13(MemoryUnit_io_csr_in_ex_tval_13),
    .io_csr_in_ex_tval_14(MemoryUnit_io_csr_in_ex_tval_14),
    .io_csr_in_ex_tval_15(MemoryUnit_io_csr_in_ex_tval_15),
    .io_csr_in_info_valid(MemoryUnit_io_csr_in_info_valid),
    .io_csr_in_info_fusel(MemoryUnit_io_csr_in_info_fusel),
    .io_csr_in_info_op(MemoryUnit_io_csr_in_info_op),
    .io_csr_in_lr_wen(MemoryUnit_io_csr_in_lr_wen),
    .io_csr_in_lr_wbit(MemoryUnit_io_csr_in_lr_wbit),
    .io_csr_in_lr_waddr(MemoryUnit_io_csr_in_lr_waddr),
    .io_csr_out_flush(MemoryUnit_io_csr_out_flush),
    .io_csr_out_target(MemoryUnit_io_csr_out_target),
    .io_csr_out_lr(MemoryUnit_io_csr_out_lr),
    .io_csr_out_lr_addr(MemoryUnit_io_csr_out_lr_addr),
    .io_writeBackStage_inst_0_pc(MemoryUnit_io_writeBackStage_inst_0_pc),
    .io_writeBackStage_inst_0_info_valid(MemoryUnit_io_writeBackStage_inst_0_info_valid),
    .io_writeBackStage_inst_0_info_fusel(MemoryUnit_io_writeBackStage_inst_0_info_fusel),
    .io_writeBackStage_inst_0_info_reg_wen(MemoryUnit_io_writeBackStage_inst_0_info_reg_wen),
    .io_writeBackStage_inst_0_info_reg_waddr(MemoryUnit_io_writeBackStage_inst_0_info_reg_waddr),
    .io_writeBackStage_inst_0_rd_info_wdata_0(MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_0),
    .io_writeBackStage_inst_0_rd_info_wdata_1(MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_1),
    .io_writeBackStage_inst_0_rd_info_wdata_2(MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_2),
    .io_writeBackStage_inst_0_rd_info_wdata_3(MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_3),
    .io_writeBackStage_inst_0_rd_info_wdata_4(MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_4),
    .io_writeBackStage_inst_0_rd_info_wdata_5(MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_5),
    .io_writeBackStage_inst_0_ex_exception_0(MemoryUnit_io_writeBackStage_inst_0_ex_exception_0),
    .io_writeBackStage_inst_0_ex_exception_1(MemoryUnit_io_writeBackStage_inst_0_ex_exception_1),
    .io_writeBackStage_inst_0_ex_exception_2(MemoryUnit_io_writeBackStage_inst_0_ex_exception_2),
    .io_writeBackStage_inst_0_ex_exception_3(MemoryUnit_io_writeBackStage_inst_0_ex_exception_3),
    .io_writeBackStage_inst_0_ex_exception_4(MemoryUnit_io_writeBackStage_inst_0_ex_exception_4),
    .io_writeBackStage_inst_0_ex_exception_5(MemoryUnit_io_writeBackStage_inst_0_ex_exception_5),
    .io_writeBackStage_inst_0_ex_exception_6(MemoryUnit_io_writeBackStage_inst_0_ex_exception_6),
    .io_writeBackStage_inst_0_ex_exception_7(MemoryUnit_io_writeBackStage_inst_0_ex_exception_7),
    .io_writeBackStage_inst_0_ex_exception_8(MemoryUnit_io_writeBackStage_inst_0_ex_exception_8),
    .io_writeBackStage_inst_0_ex_exception_9(MemoryUnit_io_writeBackStage_inst_0_ex_exception_9),
    .io_writeBackStage_inst_0_ex_exception_10(MemoryUnit_io_writeBackStage_inst_0_ex_exception_10),
    .io_writeBackStage_inst_0_ex_exception_11(MemoryUnit_io_writeBackStage_inst_0_ex_exception_11),
    .io_writeBackStage_inst_0_ex_exception_12(MemoryUnit_io_writeBackStage_inst_0_ex_exception_12),
    .io_writeBackStage_inst_0_ex_exception_13(MemoryUnit_io_writeBackStage_inst_0_ex_exception_13),
    .io_writeBackStage_inst_0_ex_exception_14(MemoryUnit_io_writeBackStage_inst_0_ex_exception_14),
    .io_writeBackStage_inst_0_ex_exception_15(MemoryUnit_io_writeBackStage_inst_0_ex_exception_15),
    .io_writeBackStage_inst_0_ex_interrupt_0(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_0),
    .io_writeBackStage_inst_0_ex_interrupt_1(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_1),
    .io_writeBackStage_inst_0_ex_interrupt_2(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_2),
    .io_writeBackStage_inst_0_ex_interrupt_3(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_3),
    .io_writeBackStage_inst_0_ex_interrupt_4(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_4),
    .io_writeBackStage_inst_0_ex_interrupt_5(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_5),
    .io_writeBackStage_inst_0_ex_interrupt_6(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_6),
    .io_writeBackStage_inst_0_ex_interrupt_7(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_7),
    .io_writeBackStage_inst_0_ex_interrupt_8(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_8),
    .io_writeBackStage_inst_0_ex_interrupt_9(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_9),
    .io_writeBackStage_inst_0_ex_interrupt_10(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_10),
    .io_writeBackStage_inst_0_ex_interrupt_11(MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_11),
    .io_writeBackStage_inst_0_ex_tval_0(MemoryUnit_io_writeBackStage_inst_0_ex_tval_0),
    .io_writeBackStage_inst_0_ex_tval_1(MemoryUnit_io_writeBackStage_inst_0_ex_tval_1),
    .io_writeBackStage_inst_0_ex_tval_2(MemoryUnit_io_writeBackStage_inst_0_ex_tval_2),
    .io_writeBackStage_inst_0_ex_tval_3(MemoryUnit_io_writeBackStage_inst_0_ex_tval_3),
    .io_writeBackStage_inst_0_ex_tval_4(MemoryUnit_io_writeBackStage_inst_0_ex_tval_4),
    .io_writeBackStage_inst_0_ex_tval_5(MemoryUnit_io_writeBackStage_inst_0_ex_tval_5),
    .io_writeBackStage_inst_0_ex_tval_6(MemoryUnit_io_writeBackStage_inst_0_ex_tval_6),
    .io_writeBackStage_inst_0_ex_tval_7(MemoryUnit_io_writeBackStage_inst_0_ex_tval_7),
    .io_writeBackStage_inst_0_ex_tval_8(MemoryUnit_io_writeBackStage_inst_0_ex_tval_8),
    .io_writeBackStage_inst_0_ex_tval_9(MemoryUnit_io_writeBackStage_inst_0_ex_tval_9),
    .io_writeBackStage_inst_0_ex_tval_10(MemoryUnit_io_writeBackStage_inst_0_ex_tval_10),
    .io_writeBackStage_inst_0_ex_tval_11(MemoryUnit_io_writeBackStage_inst_0_ex_tval_11),
    .io_writeBackStage_inst_0_ex_tval_12(MemoryUnit_io_writeBackStage_inst_0_ex_tval_12),
    .io_writeBackStage_inst_0_ex_tval_13(MemoryUnit_io_writeBackStage_inst_0_ex_tval_13),
    .io_writeBackStage_inst_0_ex_tval_14(MemoryUnit_io_writeBackStage_inst_0_ex_tval_14),
    .io_writeBackStage_inst_0_ex_tval_15(MemoryUnit_io_writeBackStage_inst_0_ex_tval_15),
    .io_writeBackStage_inst_1_pc(MemoryUnit_io_writeBackStage_inst_1_pc),
    .io_writeBackStage_inst_1_info_valid(MemoryUnit_io_writeBackStage_inst_1_info_valid),
    .io_writeBackStage_inst_1_info_fusel(MemoryUnit_io_writeBackStage_inst_1_info_fusel),
    .io_writeBackStage_inst_1_info_reg_wen(MemoryUnit_io_writeBackStage_inst_1_info_reg_wen),
    .io_writeBackStage_inst_1_info_reg_waddr(MemoryUnit_io_writeBackStage_inst_1_info_reg_waddr),
    .io_writeBackStage_inst_1_rd_info_wdata_0(MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_0),
    .io_writeBackStage_inst_1_rd_info_wdata_1(MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_1),
    .io_writeBackStage_inst_1_rd_info_wdata_2(MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_2),
    .io_writeBackStage_inst_1_rd_info_wdata_3(MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_3),
    .io_writeBackStage_inst_1_rd_info_wdata_4(MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_4),
    .io_writeBackStage_inst_1_rd_info_wdata_5(MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_5),
    .io_writeBackStage_inst_1_ex_exception_0(MemoryUnit_io_writeBackStage_inst_1_ex_exception_0),
    .io_writeBackStage_inst_1_ex_exception_1(MemoryUnit_io_writeBackStage_inst_1_ex_exception_1),
    .io_writeBackStage_inst_1_ex_exception_2(MemoryUnit_io_writeBackStage_inst_1_ex_exception_2),
    .io_writeBackStage_inst_1_ex_exception_3(MemoryUnit_io_writeBackStage_inst_1_ex_exception_3),
    .io_writeBackStage_inst_1_ex_exception_4(MemoryUnit_io_writeBackStage_inst_1_ex_exception_4),
    .io_writeBackStage_inst_1_ex_exception_5(MemoryUnit_io_writeBackStage_inst_1_ex_exception_5),
    .io_writeBackStage_inst_1_ex_exception_6(MemoryUnit_io_writeBackStage_inst_1_ex_exception_6),
    .io_writeBackStage_inst_1_ex_exception_7(MemoryUnit_io_writeBackStage_inst_1_ex_exception_7),
    .io_writeBackStage_inst_1_ex_exception_8(MemoryUnit_io_writeBackStage_inst_1_ex_exception_8),
    .io_writeBackStage_inst_1_ex_exception_9(MemoryUnit_io_writeBackStage_inst_1_ex_exception_9),
    .io_writeBackStage_inst_1_ex_exception_10(MemoryUnit_io_writeBackStage_inst_1_ex_exception_10),
    .io_writeBackStage_inst_1_ex_exception_11(MemoryUnit_io_writeBackStage_inst_1_ex_exception_11),
    .io_writeBackStage_inst_1_ex_exception_12(MemoryUnit_io_writeBackStage_inst_1_ex_exception_12),
    .io_writeBackStage_inst_1_ex_exception_13(MemoryUnit_io_writeBackStage_inst_1_ex_exception_13),
    .io_writeBackStage_inst_1_ex_exception_14(MemoryUnit_io_writeBackStage_inst_1_ex_exception_14),
    .io_writeBackStage_inst_1_ex_exception_15(MemoryUnit_io_writeBackStage_inst_1_ex_exception_15),
    .io_writeBackStage_inst_1_ex_interrupt_0(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_0),
    .io_writeBackStage_inst_1_ex_interrupt_1(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_1),
    .io_writeBackStage_inst_1_ex_interrupt_2(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_2),
    .io_writeBackStage_inst_1_ex_interrupt_3(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_3),
    .io_writeBackStage_inst_1_ex_interrupt_4(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_4),
    .io_writeBackStage_inst_1_ex_interrupt_5(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_5),
    .io_writeBackStage_inst_1_ex_interrupt_6(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_6),
    .io_writeBackStage_inst_1_ex_interrupt_7(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_7),
    .io_writeBackStage_inst_1_ex_interrupt_8(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_8),
    .io_writeBackStage_inst_1_ex_interrupt_9(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_9),
    .io_writeBackStage_inst_1_ex_interrupt_10(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_10),
    .io_writeBackStage_inst_1_ex_interrupt_11(MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_11),
    .io_writeBackStage_inst_1_ex_tval_0(MemoryUnit_io_writeBackStage_inst_1_ex_tval_0),
    .io_writeBackStage_inst_1_ex_tval_1(MemoryUnit_io_writeBackStage_inst_1_ex_tval_1),
    .io_writeBackStage_inst_1_ex_tval_2(MemoryUnit_io_writeBackStage_inst_1_ex_tval_2),
    .io_writeBackStage_inst_1_ex_tval_3(MemoryUnit_io_writeBackStage_inst_1_ex_tval_3),
    .io_writeBackStage_inst_1_ex_tval_4(MemoryUnit_io_writeBackStage_inst_1_ex_tval_4),
    .io_writeBackStage_inst_1_ex_tval_5(MemoryUnit_io_writeBackStage_inst_1_ex_tval_5),
    .io_writeBackStage_inst_1_ex_tval_6(MemoryUnit_io_writeBackStage_inst_1_ex_tval_6),
    .io_writeBackStage_inst_1_ex_tval_7(MemoryUnit_io_writeBackStage_inst_1_ex_tval_7),
    .io_writeBackStage_inst_1_ex_tval_8(MemoryUnit_io_writeBackStage_inst_1_ex_tval_8),
    .io_writeBackStage_inst_1_ex_tval_9(MemoryUnit_io_writeBackStage_inst_1_ex_tval_9),
    .io_writeBackStage_inst_1_ex_tval_10(MemoryUnit_io_writeBackStage_inst_1_ex_tval_10),
    .io_writeBackStage_inst_1_ex_tval_11(MemoryUnit_io_writeBackStage_inst_1_ex_tval_11),
    .io_writeBackStage_inst_1_ex_tval_12(MemoryUnit_io_writeBackStage_inst_1_ex_tval_12),
    .io_writeBackStage_inst_1_ex_tval_13(MemoryUnit_io_writeBackStage_inst_1_ex_tval_13),
    .io_writeBackStage_inst_1_ex_tval_14(MemoryUnit_io_writeBackStage_inst_1_ex_tval_14),
    .io_writeBackStage_inst_1_ex_tval_15(MemoryUnit_io_writeBackStage_inst_1_ex_tval_15),
    .io_dataMemory_in_access_fault(MemoryUnit_io_dataMemory_in_access_fault),
    .io_dataMemory_in_page_fault(MemoryUnit_io_dataMemory_in_page_fault),
    .io_dataMemory_in_ready(MemoryUnit_io_dataMemory_in_ready),
    .io_dataMemory_in_rdata(MemoryUnit_io_dataMemory_in_rdata),
    .io_dataMemory_out_en(MemoryUnit_io_dataMemory_out_en),
    .io_dataMemory_out_rlen(MemoryUnit_io_dataMemory_out_rlen),
    .io_dataMemory_out_wen(MemoryUnit_io_dataMemory_out_wen),
    .io_dataMemory_out_wstrb(MemoryUnit_io_dataMemory_out_wstrb),
    .io_dataMemory_out_addr(MemoryUnit_io_dataMemory_out_addr),
    .io_dataMemory_out_wdata(MemoryUnit_io_dataMemory_out_wdata)
  );
  WriteBackStage WriteBackStage ( // @[playground/src/Core.scala 36:30]
    .clock(WriteBackStage_clock),
    .reset(WriteBackStage_reset),
    .io_ctrl_allow_to_go(WriteBackStage_io_ctrl_allow_to_go),
    .io_memoryUnit_inst_0_pc(WriteBackStage_io_memoryUnit_inst_0_pc),
    .io_memoryUnit_inst_0_info_valid(WriteBackStage_io_memoryUnit_inst_0_info_valid),
    .io_memoryUnit_inst_0_info_fusel(WriteBackStage_io_memoryUnit_inst_0_info_fusel),
    .io_memoryUnit_inst_0_info_reg_wen(WriteBackStage_io_memoryUnit_inst_0_info_reg_wen),
    .io_memoryUnit_inst_0_info_reg_waddr(WriteBackStage_io_memoryUnit_inst_0_info_reg_waddr),
    .io_memoryUnit_inst_0_rd_info_wdata_0(WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_0),
    .io_memoryUnit_inst_0_rd_info_wdata_1(WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_1),
    .io_memoryUnit_inst_0_rd_info_wdata_2(WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_2),
    .io_memoryUnit_inst_0_rd_info_wdata_3(WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_3),
    .io_memoryUnit_inst_0_rd_info_wdata_5(WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_5),
    .io_memoryUnit_inst_0_ex_exception_0(WriteBackStage_io_memoryUnit_inst_0_ex_exception_0),
    .io_memoryUnit_inst_0_ex_exception_1(WriteBackStage_io_memoryUnit_inst_0_ex_exception_1),
    .io_memoryUnit_inst_0_ex_exception_2(WriteBackStage_io_memoryUnit_inst_0_ex_exception_2),
    .io_memoryUnit_inst_0_ex_exception_3(WriteBackStage_io_memoryUnit_inst_0_ex_exception_3),
    .io_memoryUnit_inst_0_ex_exception_4(WriteBackStage_io_memoryUnit_inst_0_ex_exception_4),
    .io_memoryUnit_inst_0_ex_exception_5(WriteBackStage_io_memoryUnit_inst_0_ex_exception_5),
    .io_memoryUnit_inst_0_ex_exception_6(WriteBackStage_io_memoryUnit_inst_0_ex_exception_6),
    .io_memoryUnit_inst_0_ex_exception_7(WriteBackStage_io_memoryUnit_inst_0_ex_exception_7),
    .io_memoryUnit_inst_0_ex_exception_8(WriteBackStage_io_memoryUnit_inst_0_ex_exception_8),
    .io_memoryUnit_inst_0_ex_exception_9(WriteBackStage_io_memoryUnit_inst_0_ex_exception_9),
    .io_memoryUnit_inst_0_ex_exception_11(WriteBackStage_io_memoryUnit_inst_0_ex_exception_11),
    .io_memoryUnit_inst_0_ex_exception_12(WriteBackStage_io_memoryUnit_inst_0_ex_exception_12),
    .io_memoryUnit_inst_0_ex_exception_13(WriteBackStage_io_memoryUnit_inst_0_ex_exception_13),
    .io_memoryUnit_inst_0_ex_exception_15(WriteBackStage_io_memoryUnit_inst_0_ex_exception_15),
    .io_memoryUnit_inst_0_ex_interrupt_0(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_0),
    .io_memoryUnit_inst_0_ex_interrupt_1(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_1),
    .io_memoryUnit_inst_0_ex_interrupt_2(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_2),
    .io_memoryUnit_inst_0_ex_interrupt_3(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_3),
    .io_memoryUnit_inst_0_ex_interrupt_4(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_4),
    .io_memoryUnit_inst_0_ex_interrupt_5(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_5),
    .io_memoryUnit_inst_0_ex_interrupt_6(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_6),
    .io_memoryUnit_inst_0_ex_interrupt_7(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_7),
    .io_memoryUnit_inst_0_ex_interrupt_8(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_8),
    .io_memoryUnit_inst_0_ex_interrupt_9(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_9),
    .io_memoryUnit_inst_0_ex_interrupt_10(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_10),
    .io_memoryUnit_inst_0_ex_interrupt_11(WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_11),
    .io_memoryUnit_inst_1_pc(WriteBackStage_io_memoryUnit_inst_1_pc),
    .io_memoryUnit_inst_1_info_valid(WriteBackStage_io_memoryUnit_inst_1_info_valid),
    .io_memoryUnit_inst_1_info_fusel(WriteBackStage_io_memoryUnit_inst_1_info_fusel),
    .io_memoryUnit_inst_1_info_reg_wen(WriteBackStage_io_memoryUnit_inst_1_info_reg_wen),
    .io_memoryUnit_inst_1_info_reg_waddr(WriteBackStage_io_memoryUnit_inst_1_info_reg_waddr),
    .io_memoryUnit_inst_1_rd_info_wdata_0(WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_0),
    .io_memoryUnit_inst_1_rd_info_wdata_1(WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_1),
    .io_memoryUnit_inst_1_rd_info_wdata_2(WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_2),
    .io_memoryUnit_inst_1_rd_info_wdata_3(WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_3),
    .io_memoryUnit_inst_1_rd_info_wdata_5(WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_5),
    .io_memoryUnit_inst_1_ex_exception_0(WriteBackStage_io_memoryUnit_inst_1_ex_exception_0),
    .io_memoryUnit_inst_1_ex_exception_1(WriteBackStage_io_memoryUnit_inst_1_ex_exception_1),
    .io_memoryUnit_inst_1_ex_exception_2(WriteBackStage_io_memoryUnit_inst_1_ex_exception_2),
    .io_memoryUnit_inst_1_ex_exception_3(WriteBackStage_io_memoryUnit_inst_1_ex_exception_3),
    .io_memoryUnit_inst_1_ex_exception_4(WriteBackStage_io_memoryUnit_inst_1_ex_exception_4),
    .io_memoryUnit_inst_1_ex_exception_5(WriteBackStage_io_memoryUnit_inst_1_ex_exception_5),
    .io_memoryUnit_inst_1_ex_exception_6(WriteBackStage_io_memoryUnit_inst_1_ex_exception_6),
    .io_memoryUnit_inst_1_ex_exception_7(WriteBackStage_io_memoryUnit_inst_1_ex_exception_7),
    .io_memoryUnit_inst_1_ex_exception_8(WriteBackStage_io_memoryUnit_inst_1_ex_exception_8),
    .io_memoryUnit_inst_1_ex_exception_9(WriteBackStage_io_memoryUnit_inst_1_ex_exception_9),
    .io_memoryUnit_inst_1_ex_exception_11(WriteBackStage_io_memoryUnit_inst_1_ex_exception_11),
    .io_memoryUnit_inst_1_ex_exception_12(WriteBackStage_io_memoryUnit_inst_1_ex_exception_12),
    .io_memoryUnit_inst_1_ex_exception_13(WriteBackStage_io_memoryUnit_inst_1_ex_exception_13),
    .io_memoryUnit_inst_1_ex_exception_15(WriteBackStage_io_memoryUnit_inst_1_ex_exception_15),
    .io_memoryUnit_inst_1_ex_interrupt_0(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_0),
    .io_memoryUnit_inst_1_ex_interrupt_1(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_1),
    .io_memoryUnit_inst_1_ex_interrupt_2(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_2),
    .io_memoryUnit_inst_1_ex_interrupt_3(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_3),
    .io_memoryUnit_inst_1_ex_interrupt_4(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_4),
    .io_memoryUnit_inst_1_ex_interrupt_5(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_5),
    .io_memoryUnit_inst_1_ex_interrupt_6(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_6),
    .io_memoryUnit_inst_1_ex_interrupt_7(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_7),
    .io_memoryUnit_inst_1_ex_interrupt_8(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_8),
    .io_memoryUnit_inst_1_ex_interrupt_9(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_9),
    .io_memoryUnit_inst_1_ex_interrupt_10(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_10),
    .io_memoryUnit_inst_1_ex_interrupt_11(WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_11),
    .io_writeBackUnit_inst_0_pc(WriteBackStage_io_writeBackUnit_inst_0_pc),
    .io_writeBackUnit_inst_0_info_valid(WriteBackStage_io_writeBackUnit_inst_0_info_valid),
    .io_writeBackUnit_inst_0_info_fusel(WriteBackStage_io_writeBackUnit_inst_0_info_fusel),
    .io_writeBackUnit_inst_0_info_reg_wen(WriteBackStage_io_writeBackUnit_inst_0_info_reg_wen),
    .io_writeBackUnit_inst_0_info_reg_waddr(WriteBackStage_io_writeBackUnit_inst_0_info_reg_waddr),
    .io_writeBackUnit_inst_0_rd_info_wdata_0(WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_0),
    .io_writeBackUnit_inst_0_rd_info_wdata_1(WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_1),
    .io_writeBackUnit_inst_0_rd_info_wdata_2(WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_2),
    .io_writeBackUnit_inst_0_rd_info_wdata_3(WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_3),
    .io_writeBackUnit_inst_0_rd_info_wdata_5(WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_5),
    .io_writeBackUnit_inst_0_ex_exception_0(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_0),
    .io_writeBackUnit_inst_0_ex_exception_1(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_1),
    .io_writeBackUnit_inst_0_ex_exception_2(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_2),
    .io_writeBackUnit_inst_0_ex_exception_3(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_3),
    .io_writeBackUnit_inst_0_ex_exception_4(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_4),
    .io_writeBackUnit_inst_0_ex_exception_5(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_5),
    .io_writeBackUnit_inst_0_ex_exception_6(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_6),
    .io_writeBackUnit_inst_0_ex_exception_7(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_7),
    .io_writeBackUnit_inst_0_ex_exception_8(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_8),
    .io_writeBackUnit_inst_0_ex_exception_9(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_9),
    .io_writeBackUnit_inst_0_ex_exception_11(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_11),
    .io_writeBackUnit_inst_0_ex_exception_12(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_12),
    .io_writeBackUnit_inst_0_ex_exception_13(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_13),
    .io_writeBackUnit_inst_0_ex_exception_15(WriteBackStage_io_writeBackUnit_inst_0_ex_exception_15),
    .io_writeBackUnit_inst_0_ex_interrupt_0(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_0),
    .io_writeBackUnit_inst_0_ex_interrupt_1(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_1),
    .io_writeBackUnit_inst_0_ex_interrupt_2(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_2),
    .io_writeBackUnit_inst_0_ex_interrupt_3(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_3),
    .io_writeBackUnit_inst_0_ex_interrupt_4(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_4),
    .io_writeBackUnit_inst_0_ex_interrupt_5(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_5),
    .io_writeBackUnit_inst_0_ex_interrupt_6(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_6),
    .io_writeBackUnit_inst_0_ex_interrupt_7(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_7),
    .io_writeBackUnit_inst_0_ex_interrupt_8(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_8),
    .io_writeBackUnit_inst_0_ex_interrupt_9(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_9),
    .io_writeBackUnit_inst_0_ex_interrupt_10(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_10),
    .io_writeBackUnit_inst_0_ex_interrupt_11(WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_11),
    .io_writeBackUnit_inst_1_pc(WriteBackStage_io_writeBackUnit_inst_1_pc),
    .io_writeBackUnit_inst_1_info_valid(WriteBackStage_io_writeBackUnit_inst_1_info_valid),
    .io_writeBackUnit_inst_1_info_fusel(WriteBackStage_io_writeBackUnit_inst_1_info_fusel),
    .io_writeBackUnit_inst_1_info_reg_wen(WriteBackStage_io_writeBackUnit_inst_1_info_reg_wen),
    .io_writeBackUnit_inst_1_info_reg_waddr(WriteBackStage_io_writeBackUnit_inst_1_info_reg_waddr),
    .io_writeBackUnit_inst_1_rd_info_wdata_0(WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_0),
    .io_writeBackUnit_inst_1_rd_info_wdata_1(WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_1),
    .io_writeBackUnit_inst_1_rd_info_wdata_2(WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_2),
    .io_writeBackUnit_inst_1_rd_info_wdata_3(WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_3),
    .io_writeBackUnit_inst_1_rd_info_wdata_5(WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_5),
    .io_writeBackUnit_inst_1_ex_exception_0(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_0),
    .io_writeBackUnit_inst_1_ex_exception_1(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_1),
    .io_writeBackUnit_inst_1_ex_exception_2(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_2),
    .io_writeBackUnit_inst_1_ex_exception_3(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_3),
    .io_writeBackUnit_inst_1_ex_exception_4(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_4),
    .io_writeBackUnit_inst_1_ex_exception_5(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_5),
    .io_writeBackUnit_inst_1_ex_exception_6(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_6),
    .io_writeBackUnit_inst_1_ex_exception_7(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_7),
    .io_writeBackUnit_inst_1_ex_exception_8(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_8),
    .io_writeBackUnit_inst_1_ex_exception_9(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_9),
    .io_writeBackUnit_inst_1_ex_exception_11(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_11),
    .io_writeBackUnit_inst_1_ex_exception_12(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_12),
    .io_writeBackUnit_inst_1_ex_exception_13(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_13),
    .io_writeBackUnit_inst_1_ex_exception_15(WriteBackStage_io_writeBackUnit_inst_1_ex_exception_15),
    .io_writeBackUnit_inst_1_ex_interrupt_0(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_0),
    .io_writeBackUnit_inst_1_ex_interrupt_1(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_1),
    .io_writeBackUnit_inst_1_ex_interrupt_2(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_2),
    .io_writeBackUnit_inst_1_ex_interrupt_3(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_3),
    .io_writeBackUnit_inst_1_ex_interrupt_4(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_4),
    .io_writeBackUnit_inst_1_ex_interrupt_5(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_5),
    .io_writeBackUnit_inst_1_ex_interrupt_6(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_6),
    .io_writeBackUnit_inst_1_ex_interrupt_7(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_7),
    .io_writeBackUnit_inst_1_ex_interrupt_8(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_8),
    .io_writeBackUnit_inst_1_ex_interrupt_9(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_9),
    .io_writeBackUnit_inst_1_ex_interrupt_10(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_10),
    .io_writeBackUnit_inst_1_ex_interrupt_11(WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_11)
  );
  WriteBackUnit WriteBackUnit ( // @[playground/src/Core.scala 37:30]
    .clock(WriteBackUnit_clock),
    .io_ctrl_allow_to_go(WriteBackUnit_io_ctrl_allow_to_go),
    .io_writeBackStage_inst_0_pc(WriteBackUnit_io_writeBackStage_inst_0_pc),
    .io_writeBackStage_inst_0_info_valid(WriteBackUnit_io_writeBackStage_inst_0_info_valid),
    .io_writeBackStage_inst_0_info_fusel(WriteBackUnit_io_writeBackStage_inst_0_info_fusel),
    .io_writeBackStage_inst_0_info_reg_wen(WriteBackUnit_io_writeBackStage_inst_0_info_reg_wen),
    .io_writeBackStage_inst_0_info_reg_waddr(WriteBackUnit_io_writeBackStage_inst_0_info_reg_waddr),
    .io_writeBackStage_inst_0_rd_info_wdata_0(WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_0),
    .io_writeBackStage_inst_0_rd_info_wdata_1(WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_1),
    .io_writeBackStage_inst_0_rd_info_wdata_2(WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_2),
    .io_writeBackStage_inst_0_rd_info_wdata_3(WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_3),
    .io_writeBackStage_inst_0_rd_info_wdata_5(WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_5),
    .io_writeBackStage_inst_0_ex_exception_0(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_0),
    .io_writeBackStage_inst_0_ex_exception_1(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_1),
    .io_writeBackStage_inst_0_ex_exception_2(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_2),
    .io_writeBackStage_inst_0_ex_exception_3(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_3),
    .io_writeBackStage_inst_0_ex_exception_4(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_4),
    .io_writeBackStage_inst_0_ex_exception_5(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_5),
    .io_writeBackStage_inst_0_ex_exception_6(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_6),
    .io_writeBackStage_inst_0_ex_exception_7(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_7),
    .io_writeBackStage_inst_0_ex_exception_8(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_8),
    .io_writeBackStage_inst_0_ex_exception_9(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_9),
    .io_writeBackStage_inst_0_ex_exception_11(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_11),
    .io_writeBackStage_inst_0_ex_exception_12(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_12),
    .io_writeBackStage_inst_0_ex_exception_13(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_13),
    .io_writeBackStage_inst_0_ex_exception_15(WriteBackUnit_io_writeBackStage_inst_0_ex_exception_15),
    .io_writeBackStage_inst_0_ex_interrupt_0(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_0),
    .io_writeBackStage_inst_0_ex_interrupt_1(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_1),
    .io_writeBackStage_inst_0_ex_interrupt_2(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_2),
    .io_writeBackStage_inst_0_ex_interrupt_3(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_3),
    .io_writeBackStage_inst_0_ex_interrupt_4(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_4),
    .io_writeBackStage_inst_0_ex_interrupt_5(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_5),
    .io_writeBackStage_inst_0_ex_interrupt_6(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_6),
    .io_writeBackStage_inst_0_ex_interrupt_7(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_7),
    .io_writeBackStage_inst_0_ex_interrupt_8(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_8),
    .io_writeBackStage_inst_0_ex_interrupt_9(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_9),
    .io_writeBackStage_inst_0_ex_interrupt_10(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_10),
    .io_writeBackStage_inst_0_ex_interrupt_11(WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_11),
    .io_writeBackStage_inst_1_pc(WriteBackUnit_io_writeBackStage_inst_1_pc),
    .io_writeBackStage_inst_1_info_valid(WriteBackUnit_io_writeBackStage_inst_1_info_valid),
    .io_writeBackStage_inst_1_info_fusel(WriteBackUnit_io_writeBackStage_inst_1_info_fusel),
    .io_writeBackStage_inst_1_info_reg_wen(WriteBackUnit_io_writeBackStage_inst_1_info_reg_wen),
    .io_writeBackStage_inst_1_info_reg_waddr(WriteBackUnit_io_writeBackStage_inst_1_info_reg_waddr),
    .io_writeBackStage_inst_1_rd_info_wdata_0(WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_0),
    .io_writeBackStage_inst_1_rd_info_wdata_1(WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_1),
    .io_writeBackStage_inst_1_rd_info_wdata_2(WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_2),
    .io_writeBackStage_inst_1_rd_info_wdata_3(WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_3),
    .io_writeBackStage_inst_1_rd_info_wdata_5(WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_5),
    .io_writeBackStage_inst_1_ex_exception_0(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_0),
    .io_writeBackStage_inst_1_ex_exception_1(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_1),
    .io_writeBackStage_inst_1_ex_exception_2(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_2),
    .io_writeBackStage_inst_1_ex_exception_3(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_3),
    .io_writeBackStage_inst_1_ex_exception_4(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_4),
    .io_writeBackStage_inst_1_ex_exception_5(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_5),
    .io_writeBackStage_inst_1_ex_exception_6(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_6),
    .io_writeBackStage_inst_1_ex_exception_7(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_7),
    .io_writeBackStage_inst_1_ex_exception_8(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_8),
    .io_writeBackStage_inst_1_ex_exception_9(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_9),
    .io_writeBackStage_inst_1_ex_exception_11(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_11),
    .io_writeBackStage_inst_1_ex_exception_12(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_12),
    .io_writeBackStage_inst_1_ex_exception_13(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_13),
    .io_writeBackStage_inst_1_ex_exception_15(WriteBackUnit_io_writeBackStage_inst_1_ex_exception_15),
    .io_writeBackStage_inst_1_ex_interrupt_0(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_0),
    .io_writeBackStage_inst_1_ex_interrupt_1(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_1),
    .io_writeBackStage_inst_1_ex_interrupt_2(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_2),
    .io_writeBackStage_inst_1_ex_interrupt_3(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_3),
    .io_writeBackStage_inst_1_ex_interrupt_4(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_4),
    .io_writeBackStage_inst_1_ex_interrupt_5(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_5),
    .io_writeBackStage_inst_1_ex_interrupt_6(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_6),
    .io_writeBackStage_inst_1_ex_interrupt_7(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_7),
    .io_writeBackStage_inst_1_ex_interrupt_8(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_8),
    .io_writeBackStage_inst_1_ex_interrupt_9(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_9),
    .io_writeBackStage_inst_1_ex_interrupt_10(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_10),
    .io_writeBackStage_inst_1_ex_interrupt_11(WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_11),
    .io_regfile_0_wen(WriteBackUnit_io_regfile_0_wen),
    .io_regfile_0_waddr(WriteBackUnit_io_regfile_0_waddr),
    .io_regfile_0_wdata(WriteBackUnit_io_regfile_0_wdata),
    .io_regfile_1_wen(WriteBackUnit_io_regfile_1_wen),
    .io_regfile_1_waddr(WriteBackUnit_io_regfile_1_waddr),
    .io_regfile_1_wdata(WriteBackUnit_io_regfile_1_wdata),
    .io_debug_wb_pc(WriteBackUnit_io_debug_wb_pc),
    .io_debug_wb_rf_wen(WriteBackUnit_io_debug_wb_rf_wen),
    .io_debug_wb_rf_wnum(WriteBackUnit_io_debug_wb_rf_wnum),
    .io_debug_wb_rf_wdata(WriteBackUnit_io_debug_wb_rf_wdata)
  );
  Tlb Tlb ( // @[playground/src/Core.scala 38:30]
    .clock(Tlb_clock),
    .reset(Tlb_reset),
    .io_icache_en(Tlb_io_icache_en),
    .io_icache_vaddr(Tlb_io_icache_vaddr),
    .io_icache_complete_single_request(Tlb_io_icache_complete_single_request),
    .io_icache_uncached(Tlb_io_icache_uncached),
    .io_icache_hit(Tlb_io_icache_hit),
    .io_icache_ptag(Tlb_io_icache_ptag),
    .io_icache_paddr(Tlb_io_icache_paddr),
    .io_icache_page_fault(Tlb_io_icache_page_fault),
    .io_dcache_en(Tlb_io_dcache_en),
    .io_dcache_vaddr(Tlb_io_dcache_vaddr),
    .io_dcache_complete_single_request(Tlb_io_dcache_complete_single_request),
    .io_dcache_uncached(Tlb_io_dcache_uncached),
    .io_dcache_hit(Tlb_io_dcache_hit),
    .io_dcache_ptag(Tlb_io_dcache_ptag),
    .io_dcache_paddr(Tlb_io_dcache_paddr),
    .io_dcache_page_fault(Tlb_io_dcache_page_fault),
    .io_dcache_access_type(Tlb_io_dcache_access_type),
    .io_dcache_ptw_vpn_ready(Tlb_io_dcache_ptw_vpn_ready),
    .io_dcache_ptw_vpn_valid(Tlb_io_dcache_ptw_vpn_valid),
    .io_dcache_ptw_vpn_bits(Tlb_io_dcache_ptw_vpn_bits),
    .io_dcache_ptw_access_type(Tlb_io_dcache_ptw_access_type),
    .io_dcache_ptw_pte_valid(Tlb_io_dcache_ptw_pte_valid),
    .io_dcache_ptw_pte_bits_page_fault(Tlb_io_dcache_ptw_pte_bits_page_fault),
    .io_dcache_ptw_pte_bits_entry_ppn(Tlb_io_dcache_ptw_pte_bits_entry_ppn),
    .io_dcache_ptw_pte_bits_entry_flag_d(Tlb_io_dcache_ptw_pte_bits_entry_flag_d),
    .io_dcache_ptw_pte_bits_entry_flag_g(Tlb_io_dcache_ptw_pte_bits_entry_flag_g),
    .io_dcache_ptw_pte_bits_entry_flag_u(Tlb_io_dcache_ptw_pte_bits_entry_flag_u),
    .io_dcache_ptw_pte_bits_entry_flag_x(Tlb_io_dcache_ptw_pte_bits_entry_flag_x),
    .io_dcache_ptw_pte_bits_entry_flag_w(Tlb_io_dcache_ptw_pte_bits_entry_flag_w),
    .io_dcache_ptw_pte_bits_entry_flag_r(Tlb_io_dcache_ptw_pte_bits_entry_flag_r),
    .io_dcache_ptw_pte_bits_entry_flag_v(Tlb_io_dcache_ptw_pte_bits_entry_flag_v),
    .io_dcache_ptw_pte_bits_rmask(Tlb_io_dcache_ptw_pte_bits_rmask),
    .io_dcache_csr_satp(Tlb_io_dcache_csr_satp),
    .io_dcache_csr_mstatus(Tlb_io_dcache_csr_mstatus),
    .io_dcache_csr_imode(Tlb_io_dcache_csr_imode),
    .io_dcache_csr_dmode(Tlb_io_dcache_csr_dmode),
    .io_csr_satp(Tlb_io_csr_satp),
    .io_csr_mstatus(Tlb_io_csr_mstatus),
    .io_csr_imode(Tlb_io_csr_imode),
    .io_csr_dmode(Tlb_io_csr_dmode),
    .io_sfence_vma_valid(Tlb_io_sfence_vma_valid),
    .io_sfence_vma_src_info_src1_data(Tlb_io_sfence_vma_src_info_src1_data),
    .io_sfence_vma_src_info_src2_data(Tlb_io_sfence_vma_src_info_src2_data)
  );
  assign io_inst_req = ~InstFifo_io_full & ~reset; // @[playground/src/Core.scala 136:33]
  assign io_inst_complete_single_request = Ctrl_io_fetchUnit_allow_to_go; // @[playground/src/Core.scala 138:35]
  assign io_inst_addr_0 = FetchUnit_io_iCache_pc; // @[playground/src/Core.scala 56:31]
  assign io_inst_addr_1 = FetchUnit_io_iCache_pc_next; // @[playground/src/Core.scala 57:31]
  assign io_inst_fence_i = MemoryUnit_io_ctrl_fence_i; // @[playground/src/Core.scala 132:24]
  assign io_inst_dcache_stall = ~io_data_dcache_ready; // @[playground/src/Core.scala 134:27]
  assign io_inst_tlb_uncached = Tlb_io_icache_uncached; // @[playground/src/Core.scala 40:14]
  assign io_inst_tlb_hit = Tlb_io_icache_hit; // @[playground/src/Core.scala 40:14]
  assign io_inst_tlb_ptag = Tlb_io_icache_ptag; // @[playground/src/Core.scala 40:14]
  assign io_inst_tlb_paddr = Tlb_io_icache_paddr; // @[playground/src/Core.scala 40:14]
  assign io_inst_tlb_page_fault = Tlb_io_icache_page_fault; // @[playground/src/Core.scala 40:14]
  assign io_data_exe_addr = ExecuteUnit_io_dataMemory_addr; // @[playground/src/Core.scala 119:41]
  assign io_data_addr = MemoryUnit_io_dataMemory_out_addr; // @[playground/src/Core.scala 117:41]
  assign io_data_rlen = MemoryUnit_io_dataMemory_out_rlen; // @[playground/src/Core.scala 114:41]
  assign io_data_en = MemoryUnit_io_dataMemory_out_en; // @[playground/src/Core.scala 113:41]
  assign io_data_wen = MemoryUnit_io_dataMemory_out_wen; // @[playground/src/Core.scala 115:41]
  assign io_data_wdata = MemoryUnit_io_dataMemory_out_wdata; // @[playground/src/Core.scala 116:41]
  assign io_data_complete_single_request = Ctrl_io_memoryUnit_allow_to_go | Ctrl_io_memoryUnit_complete_single_request; // @[playground/src/Core.scala 139:66]
  assign io_data_fence_i = MemoryUnit_io_ctrl_fence_i; // @[playground/src/Core.scala 133:24]
  assign io_data_wstrb = MemoryUnit_io_dataMemory_out_wstrb; // @[playground/src/Core.scala 118:41]
  assign io_data_tlb_uncached = Tlb_io_dcache_uncached; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_hit = Tlb_io_dcache_hit; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_ptag = Tlb_io_dcache_ptag; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_paddr = Tlb_io_dcache_paddr; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_page_fault = Tlb_io_dcache_page_fault; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_ptw_vpn_valid = Tlb_io_dcache_ptw_vpn_valid; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_ptw_vpn_bits = Tlb_io_dcache_ptw_vpn_bits; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_ptw_access_type = Tlb_io_dcache_ptw_access_type; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_csr_satp = Tlb_io_dcache_csr_satp; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_csr_mstatus = Tlb_io_dcache_csr_mstatus; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_csr_imode = Tlb_io_dcache_csr_imode; // @[playground/src/Core.scala 41:14]
  assign io_data_tlb_csr_dmode = Tlb_io_dcache_csr_dmode; // @[playground/src/Core.scala 41:14]
  assign io_debug_wb_pc = WriteBackUnit_io_debug_wb_pc; // @[playground/src/Core.scala 129:12]
  assign io_debug_wb_rf_wen = WriteBackUnit_io_debug_wb_rf_wen; // @[playground/src/Core.scala 129:12]
  assign io_debug_wb_rf_wnum = WriteBackUnit_io_debug_wb_rf_wnum; // @[playground/src/Core.scala 129:12]
  assign io_debug_wb_rf_wdata = WriteBackUnit_io_debug_wb_rf_wdata; // @[playground/src/Core.scala 129:12]
  assign Ctrl_io_cacheCtrl_iCache_stall = io_inst_icache_stall; // @[playground/src/Core.scala 49:31]
  assign Ctrl_io_decodeUnit_inst0_src1_ren = DecodeUnit_io_ctrl_inst0_src1_ren; // @[playground/src/Core.scala 45:19]
  assign Ctrl_io_decodeUnit_inst0_src1_raddr = DecodeUnit_io_ctrl_inst0_src1_raddr; // @[playground/src/Core.scala 45:19]
  assign Ctrl_io_decodeUnit_inst0_src2_ren = DecodeUnit_io_ctrl_inst0_src2_ren; // @[playground/src/Core.scala 45:19]
  assign Ctrl_io_decodeUnit_inst0_src2_raddr = DecodeUnit_io_ctrl_inst0_src2_raddr; // @[playground/src/Core.scala 45:19]
  assign Ctrl_io_decodeUnit_branch = DecodeUnit_io_ctrl_branch; // @[playground/src/Core.scala 45:19]
  assign Ctrl_io_executeUnit_inst_0_is_load = ExecuteUnit_io_ctrl_inst_0_is_load; // @[playground/src/Core.scala 46:20]
  assign Ctrl_io_executeUnit_inst_0_reg_waddr = ExecuteUnit_io_ctrl_inst_0_reg_waddr; // @[playground/src/Core.scala 46:20]
  assign Ctrl_io_executeUnit_inst_1_is_load = ExecuteUnit_io_ctrl_inst_1_is_load; // @[playground/src/Core.scala 46:20]
  assign Ctrl_io_executeUnit_inst_1_reg_waddr = ExecuteUnit_io_ctrl_inst_1_reg_waddr; // @[playground/src/Core.scala 46:20]
  assign Ctrl_io_executeUnit_flush = ExecuteUnit_io_ctrl_flush; // @[playground/src/Core.scala 46:20]
  assign Ctrl_io_executeUnit_fu_stall = ExecuteUnit_io_ctrl_fu_stall; // @[playground/src/Core.scala 46:20]
  assign Ctrl_io_memoryUnit_flush = MemoryUnit_io_ctrl_flush; // @[playground/src/Core.scala 47:19]
  assign Ctrl_io_memoryUnit_mem_stall = MemoryUnit_io_ctrl_mem_stall; // @[playground/src/Core.scala 47:19]
  assign Ctrl_io_memoryUnit_complete_single_request = MemoryUnit_io_ctrl_complete_single_request; // @[playground/src/Core.scala 47:19]
  assign FetchUnit_clock = clock;
  assign FetchUnit_reset = reset;
  assign FetchUnit_io_memory_flush = MemoryUnit_io_fetchUnit_flush; // @[playground/src/Core.scala 51:20]
  assign FetchUnit_io_memory_target = MemoryUnit_io_fetchUnit_target; // @[playground/src/Core.scala 51:20]
  assign FetchUnit_io_decode_branch = DecodeUnit_io_fetchUnit_branch; // @[playground/src/Core.scala 53:20]
  assign FetchUnit_io_decode_target = DecodeUnit_io_fetchUnit_target; // @[playground/src/Core.scala 53:20]
  assign FetchUnit_io_execute_flush = ExecuteUnit_io_fetchUnit_flush; // @[playground/src/Core.scala 52:21]
  assign FetchUnit_io_execute_target = ExecuteUnit_io_fetchUnit_target; // @[playground/src/Core.scala 52:21]
  assign FetchUnit_io_instFifo_full = InstFifo_io_full; // @[playground/src/Core.scala 54:31]
  assign FetchUnit_io_iCache_inst_valid_0 = io_inst_inst_valid_0; // @[playground/src/Core.scala 55:31]
  assign FetchUnit_io_iCache_inst_valid_1 = io_inst_inst_valid_1; // @[playground/src/Core.scala 55:31]
  assign BranchPredictorUnit_clock = clock;
  assign BranchPredictorUnit_reset = reset;
  assign BranchPredictorUnit_io_decode_pc = DecodeUnit_io_bpu_pc; // @[playground/src/Core.scala 62:14]
  assign BranchPredictorUnit_io_decode_info_valid = DecodeUnit_io_bpu_info_valid; // @[playground/src/Core.scala 62:14]
  assign BranchPredictorUnit_io_decode_info_fusel = DecodeUnit_io_bpu_info_fusel; // @[playground/src/Core.scala 62:14]
  assign BranchPredictorUnit_io_decode_info_op = DecodeUnit_io_bpu_info_op; // @[playground/src/Core.scala 62:14]
  assign BranchPredictorUnit_io_decode_info_imm = DecodeUnit_io_bpu_info_imm; // @[playground/src/Core.scala 62:14]
  assign BranchPredictorUnit_io_decode_pht_index = DecodeUnit_io_bpu_pht_index; // @[playground/src/Core.scala 62:14]
  assign BranchPredictorUnit_io_instBuffer_pc_0 = InstFifo_io_write_0_pc; // @[playground/src/Core.scala 70:39]
  assign BranchPredictorUnit_io_instBuffer_pc_1 = InstFifo_io_write_1_pc; // @[playground/src/Core.scala 70:39]
  assign BranchPredictorUnit_io_execute_pc = ExecuteUnit_io_bpu_pc; // @[playground/src/Core.scala 63:15]
  assign BranchPredictorUnit_io_execute_update_pht_index = ExecuteUnit_io_bpu_update_pht_index; // @[playground/src/Core.scala 63:15]
  assign BranchPredictorUnit_io_execute_branch_inst = ExecuteUnit_io_bpu_branch_inst; // @[playground/src/Core.scala 63:15]
  assign BranchPredictorUnit_io_execute_branch = ExecuteUnit_io_bpu_branch; // @[playground/src/Core.scala 63:15]
  assign InstFifo_clock = clock;
  assign InstFifo_reset = reset;
  assign InstFifo_io_do_flush = Ctrl_io_decodeUnit_do_flush; // @[playground/src/Core.scala 65:21]
  assign InstFifo_io_wen_0 = io_inst_inst_valid_0; // @[playground/src/Core.scala 71:39]
  assign InstFifo_io_wen_1 = io_inst_inst_valid_1; // @[playground/src/Core.scala 71:39]
  assign InstFifo_io_write_0_inst = io_inst_inst_0; // @[playground/src/Core.scala 73:39]
  assign InstFifo_io_write_0_pht_index = BranchPredictorUnit_io_instBuffer_pht_index_0; // @[playground/src/Core.scala 69:39]
  assign InstFifo_io_write_0_addr_misaligned = io_inst_addr_misaligned; // @[playground/src/Core.scala 76:39]
  assign InstFifo_io_write_0_access_fault = io_inst_access_fault; // @[playground/src/Core.scala 74:39]
  assign InstFifo_io_write_0_page_fault = io_inst_page_fault; // @[playground/src/Core.scala 75:39]
  assign InstFifo_io_write_0_pc = _T[63:0]; // @[playground/src/Core.scala 72:58]
  assign InstFifo_io_write_1_inst = io_inst_inst_1; // @[playground/src/Core.scala 73:39]
  assign InstFifo_io_write_1_pht_index = BranchPredictorUnit_io_instBuffer_pht_index_1; // @[playground/src/Core.scala 69:39]
  assign InstFifo_io_write_1_addr_misaligned = io_inst_addr_misaligned; // @[playground/src/Core.scala 76:39]
  assign InstFifo_io_write_1_access_fault = io_inst_access_fault; // @[playground/src/Core.scala 74:39]
  assign InstFifo_io_write_1_page_fault = io_inst_page_fault; // @[playground/src/Core.scala 75:39]
  assign InstFifo_io_write_1_pc = io_inst_addr_0 + 64'h4; // @[playground/src/Core.scala 72:58]
  assign InstFifo_io_decoderUint_allow_to_go_0 = DecodeUnit_io_instFifo_allow_to_go_0; // @[playground/src/Core.scala 66:24]
  assign InstFifo_io_decoderUint_allow_to_go_1 = DecodeUnit_io_instFifo_allow_to_go_1; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_0_inst = InstFifo_io_decoderUint_inst_0_inst; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_0_pht_index = InstFifo_io_decoderUint_inst_0_pht_index; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_0_addr_misaligned = InstFifo_io_decoderUint_inst_0_addr_misaligned; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_0_access_fault = InstFifo_io_decoderUint_inst_0_access_fault; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_0_page_fault = InstFifo_io_decoderUint_inst_0_page_fault; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_0_pc = InstFifo_io_decoderUint_inst_0_pc; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_1_inst = InstFifo_io_decoderUint_inst_1_inst; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_1_addr_misaligned = InstFifo_io_decoderUint_inst_1_addr_misaligned; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_1_access_fault = InstFifo_io_decoderUint_inst_1_access_fault; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_1_page_fault = InstFifo_io_decoderUint_inst_1_page_fault; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_inst_1_pc = InstFifo_io_decoderUint_inst_1_pc; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_info_empty = InstFifo_io_decoderUint_info_empty; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_instFifo_info_almost_empty = InstFifo_io_decoderUint_info_almost_empty; // @[playground/src/Core.scala 66:24]
  assign DecodeUnit_io_regfile_0_src1_rdata = ARegFile_io_read_0_src1_rdata; // @[playground/src/Core.scala 79:22]
  assign DecodeUnit_io_regfile_0_src2_rdata = ARegFile_io_read_0_src2_rdata; // @[playground/src/Core.scala 79:22]
  assign DecodeUnit_io_regfile_1_src1_rdata = ARegFile_io_read_1_src1_rdata; // @[playground/src/Core.scala 79:22]
  assign DecodeUnit_io_regfile_1_src2_rdata = ARegFile_io_read_1_src2_rdata; // @[playground/src/Core.scala 79:22]
  assign DecodeUnit_io_forward_0_exe_wen = ExecuteUnit_io_decodeUnit_forward_0_exe_wen; // @[playground/src/Core.scala 81:35]
  assign DecodeUnit_io_forward_0_exe_waddr = ExecuteUnit_io_decodeUnit_forward_0_exe_waddr; // @[playground/src/Core.scala 81:35]
  assign DecodeUnit_io_forward_0_exe_wdata = ExecuteUnit_io_decodeUnit_forward_0_exe_wdata; // @[playground/src/Core.scala 81:35]
  assign DecodeUnit_io_forward_0_is_load = ExecuteUnit_io_decodeUnit_forward_0_is_load; // @[playground/src/Core.scala 82:35]
  assign DecodeUnit_io_forward_0_mem_wen = MemoryUnit_io_decodeUnit_0_wen; // @[playground/src/Core.scala 83:35]
  assign DecodeUnit_io_forward_0_mem_waddr = MemoryUnit_io_decodeUnit_0_waddr; // @[playground/src/Core.scala 83:35]
  assign DecodeUnit_io_forward_0_mem_wdata = MemoryUnit_io_decodeUnit_0_wdata; // @[playground/src/Core.scala 83:35]
  assign DecodeUnit_io_forward_1_exe_wen = ExecuteUnit_io_decodeUnit_forward_1_exe_wen; // @[playground/src/Core.scala 81:35]
  assign DecodeUnit_io_forward_1_exe_waddr = ExecuteUnit_io_decodeUnit_forward_1_exe_waddr; // @[playground/src/Core.scala 81:35]
  assign DecodeUnit_io_forward_1_exe_wdata = ExecuteUnit_io_decodeUnit_forward_1_exe_wdata; // @[playground/src/Core.scala 81:35]
  assign DecodeUnit_io_forward_1_is_load = ExecuteUnit_io_decodeUnit_forward_1_is_load; // @[playground/src/Core.scala 82:35]
  assign DecodeUnit_io_forward_1_mem_wen = MemoryUnit_io_decodeUnit_1_wen; // @[playground/src/Core.scala 83:35]
  assign DecodeUnit_io_forward_1_mem_waddr = MemoryUnit_io_decodeUnit_1_waddr; // @[playground/src/Core.scala 83:35]
  assign DecodeUnit_io_forward_1_mem_wdata = MemoryUnit_io_decodeUnit_1_wdata; // @[playground/src/Core.scala 83:35]
  assign DecodeUnit_io_csr_mode = Csr_io_decodeUnit_mode; // @[playground/src/Core.scala 85:18]
  assign DecodeUnit_io_csr_interrupt = Csr_io_decodeUnit_interrupt; // @[playground/src/Core.scala 85:18]
  assign DecodeUnit_io_bpu_branch_inst = BranchPredictorUnit_io_decode_branch_inst; // @[playground/src/Core.scala 62:14]
  assign DecodeUnit_io_bpu_branch = BranchPredictorUnit_io_decode_branch; // @[playground/src/Core.scala 62:14]
  assign DecodeUnit_io_bpu_target = BranchPredictorUnit_io_decode_target; // @[playground/src/Core.scala 62:14]
  assign DecodeUnit_io_bpu_update_pht_index = BranchPredictorUnit_io_decode_update_pht_index; // @[playground/src/Core.scala 62:14]
  assign DecodeUnit_io_ctrl_allow_to_go = Ctrl_io_decodeUnit_allow_to_go; // @[playground/src/Core.scala 45:19]
  assign ARegFile_clock = clock;
  assign ARegFile_reset = reset;
  assign ARegFile_io_read_0_src1_raddr = DecodeUnit_io_regfile_0_src1_raddr; // @[playground/src/Core.scala 79:22]
  assign ARegFile_io_read_0_src2_raddr = DecodeUnit_io_regfile_0_src2_raddr; // @[playground/src/Core.scala 79:22]
  assign ARegFile_io_read_1_src1_raddr = DecodeUnit_io_regfile_1_src1_raddr; // @[playground/src/Core.scala 79:22]
  assign ARegFile_io_read_1_src2_raddr = DecodeUnit_io_regfile_1_src2_raddr; // @[playground/src/Core.scala 79:22]
  assign ARegFile_io_write_0_wen = WriteBackUnit_io_regfile_0_wen; // @[playground/src/Core.scala 127:17]
  assign ARegFile_io_write_0_waddr = WriteBackUnit_io_regfile_0_waddr; // @[playground/src/Core.scala 127:17]
  assign ARegFile_io_write_0_wdata = WriteBackUnit_io_regfile_0_wdata; // @[playground/src/Core.scala 127:17]
  assign ARegFile_io_write_1_wen = WriteBackUnit_io_regfile_1_wen; // @[playground/src/Core.scala 127:17]
  assign ARegFile_io_write_1_waddr = WriteBackUnit_io_regfile_1_waddr; // @[playground/src/Core.scala 127:17]
  assign ARegFile_io_write_1_wdata = WriteBackUnit_io_regfile_1_wdata; // @[playground/src/Core.scala 127:17]
  assign ExecuteStage_clock = clock;
  assign ExecuteStage_reset = reset;
  assign ExecuteStage_io_ctrl_allow_to_go_0 = DecodeUnit_io_instFifo_allow_to_go_0; // @[playground/src/Core.scala 94:38]
  assign ExecuteStage_io_ctrl_allow_to_go_1 = DecodeUnit_io_instFifo_allow_to_go_1; // @[playground/src/Core.scala 94:38]
  assign ExecuteStage_io_ctrl_clear_0 = Ctrl_io_memoryUnit_do_flush | Ctrl_io_executeUnit_do_flush | _T_6; // @[playground/src/Core.scala 91:61]
  assign ExecuteStage_io_ctrl_clear_1 = Ctrl_io_memoryUnit_do_flush | Ctrl_io_executeUnit_do_flush | _T_10; // @[playground/src/Core.scala 91:61]
  assign ExecuteStage_io_decodeUnit_inst_0_pc = DecodeUnit_io_executeStage_inst_0_pc; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_valid = DecodeUnit_io_executeStage_inst_0_info_valid; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_fusel = DecodeUnit_io_executeStage_inst_0_info_fusel; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_op = DecodeUnit_io_executeStage_inst_0_info_op; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_reg_wen = DecodeUnit_io_executeStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_reg_waddr = DecodeUnit_io_executeStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_imm = DecodeUnit_io_executeStage_inst_0_info_imm; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_info_inst = DecodeUnit_io_executeStage_inst_0_info_inst; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_src_info_src1_data = DecodeUnit_io_executeStage_inst_0_src_info_src1_data; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_src_info_src2_data = DecodeUnit_io_executeStage_inst_0_src_info_src2_data; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_0 = DecodeUnit_io_executeStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_1 = DecodeUnit_io_executeStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_2 = DecodeUnit_io_executeStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_3 = DecodeUnit_io_executeStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_8 = DecodeUnit_io_executeStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_9 = DecodeUnit_io_executeStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_11 = DecodeUnit_io_executeStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_exception_12 = DecodeUnit_io_executeStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_0 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_1 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_2 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_3 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_4 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_5 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_6 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_7 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_8 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_9 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_10 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_interrupt_11 = DecodeUnit_io_executeStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_tval_0 = DecodeUnit_io_executeStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_tval_1 = DecodeUnit_io_executeStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_tval_2 = DecodeUnit_io_executeStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_0_ex_tval_12 = DecodeUnit_io_executeStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_pc = DecodeUnit_io_executeStage_inst_1_pc; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_valid = DecodeUnit_io_executeStage_inst_1_info_valid; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_fusel = DecodeUnit_io_executeStage_inst_1_info_fusel; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_op = DecodeUnit_io_executeStage_inst_1_info_op; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_reg_wen = DecodeUnit_io_executeStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_reg_waddr = DecodeUnit_io_executeStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_imm = DecodeUnit_io_executeStage_inst_1_info_imm; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_info_inst = DecodeUnit_io_executeStage_inst_1_info_inst; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_src_info_src1_data = DecodeUnit_io_executeStage_inst_1_src_info_src1_data; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_src_info_src2_data = DecodeUnit_io_executeStage_inst_1_src_info_src2_data; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_0 = DecodeUnit_io_executeStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_1 = DecodeUnit_io_executeStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_2 = DecodeUnit_io_executeStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_3 = DecodeUnit_io_executeStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_8 = DecodeUnit_io_executeStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_9 = DecodeUnit_io_executeStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_11 = DecodeUnit_io_executeStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_exception_12 = DecodeUnit_io_executeStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_0 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_1 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_2 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_3 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_4 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_5 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_6 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_7 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_8 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_9 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_10 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_interrupt_11 = DecodeUnit_io_executeStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_tval_0 = DecodeUnit_io_executeStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_tval_1 = DecodeUnit_io_executeStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_tval_2 = DecodeUnit_io_executeStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_inst_1_ex_tval_12 = DecodeUnit_io_executeStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_jump_branch_info_jump_regiser =
    DecodeUnit_io_executeStage_jump_branch_info_jump_regiser; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_jump_branch_info_branch_inst =
    DecodeUnit_io_executeStage_jump_branch_info_branch_inst; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_jump_branch_info_pred_branch =
    DecodeUnit_io_executeStage_jump_branch_info_pred_branch; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_jump_branch_info_branch_target =
    DecodeUnit_io_executeStage_jump_branch_info_branch_target; // @[playground/src/Core.scala 86:27]
  assign ExecuteStage_io_decodeUnit_jump_branch_info_update_pht_index =
    DecodeUnit_io_executeStage_jump_branch_info_update_pht_index; // @[playground/src/Core.scala 86:27]
  assign ExecuteUnit_clock = clock;
  assign ExecuteUnit_reset = reset;
  assign ExecuteUnit_io_ctrl_allow_to_go = Ctrl_io_executeUnit_allow_to_go; // @[playground/src/Core.scala 46:20]
  assign ExecuteUnit_io_ctrl_fu_allow_to_go = Ctrl_io_executeUnit_fu_allow_to_go; // @[playground/src/Core.scala 46:20]
  assign ExecuteUnit_io_executeStage_inst_0_pc = ExecuteStage_io_executeUnit_inst_0_pc; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_valid = ExecuteStage_io_executeUnit_inst_0_info_valid; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_fusel = ExecuteStage_io_executeUnit_inst_0_info_fusel; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_op = ExecuteStage_io_executeUnit_inst_0_info_op; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_reg_wen = ExecuteStage_io_executeUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_reg_waddr = ExecuteStage_io_executeUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_imm = ExecuteStage_io_executeUnit_inst_0_info_imm; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_info_inst = ExecuteStage_io_executeUnit_inst_0_info_inst; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_src_info_src1_data = ExecuteStage_io_executeUnit_inst_0_src_info_src1_data; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_src_info_src2_data = ExecuteStage_io_executeUnit_inst_0_src_info_src2_data; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_0 = ExecuteStage_io_executeUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_1 = ExecuteStage_io_executeUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_2 = ExecuteStage_io_executeUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_3 = ExecuteStage_io_executeUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_8 = ExecuteStage_io_executeUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_9 = ExecuteStage_io_executeUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_11 = ExecuteStage_io_executeUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_exception_12 = ExecuteStage_io_executeUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_0 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_1 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_2 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_3 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_4 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_5 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_6 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_7 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_8 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_9 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_10 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_interrupt_11 = ExecuteStage_io_executeUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_tval_0 = ExecuteStage_io_executeUnit_inst_0_ex_tval_0; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_tval_1 = ExecuteStage_io_executeUnit_inst_0_ex_tval_1; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_tval_2 = ExecuteStage_io_executeUnit_inst_0_ex_tval_2; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_0_ex_tval_12 = ExecuteStage_io_executeUnit_inst_0_ex_tval_12; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_pc = ExecuteStage_io_executeUnit_inst_1_pc; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_valid = ExecuteStage_io_executeUnit_inst_1_info_valid; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_fusel = ExecuteStage_io_executeUnit_inst_1_info_fusel; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_op = ExecuteStage_io_executeUnit_inst_1_info_op; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_reg_wen = ExecuteStage_io_executeUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_reg_waddr = ExecuteStage_io_executeUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_imm = ExecuteStage_io_executeUnit_inst_1_info_imm; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_info_inst = ExecuteStage_io_executeUnit_inst_1_info_inst; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_src_info_src1_data = ExecuteStage_io_executeUnit_inst_1_src_info_src1_data; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_src_info_src2_data = ExecuteStage_io_executeUnit_inst_1_src_info_src2_data; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_0 = ExecuteStage_io_executeUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_1 = ExecuteStage_io_executeUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_2 = ExecuteStage_io_executeUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_3 = ExecuteStage_io_executeUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_8 = ExecuteStage_io_executeUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_9 = ExecuteStage_io_executeUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_11 = ExecuteStage_io_executeUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_exception_12 = ExecuteStage_io_executeUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_0 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_1 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_2 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_3 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_4 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_5 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_6 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_7 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_8 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_9 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_10 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_interrupt_11 = ExecuteStage_io_executeUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_tval_0 = ExecuteStage_io_executeUnit_inst_1_ex_tval_0; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_tval_1 = ExecuteStage_io_executeUnit_inst_1_ex_tval_1; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_tval_2 = ExecuteStage_io_executeUnit_inst_1_ex_tval_2; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_inst_1_ex_tval_12 = ExecuteStage_io_executeUnit_inst_1_ex_tval_12; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_jump_branch_info_jump_regiser =
    ExecuteStage_io_executeUnit_jump_branch_info_jump_regiser; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_jump_branch_info_branch_inst =
    ExecuteStage_io_executeUnit_jump_branch_info_branch_inst; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_jump_branch_info_pred_branch =
    ExecuteStage_io_executeUnit_jump_branch_info_pred_branch; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_jump_branch_info_branch_target =
    ExecuteStage_io_executeUnit_jump_branch_info_branch_target; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_executeStage_jump_branch_info_update_pht_index =
    ExecuteStage_io_executeUnit_jump_branch_info_update_pht_index; // @[playground/src/Core.scala 96:28]
  assign ExecuteUnit_io_csr_out_rdata = Csr_io_executeUnit_out_rdata; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_1 = Csr_io_executeUnit_out_ex_exception_1; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_2 = Csr_io_executeUnit_out_ex_exception_2; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_3 = Csr_io_executeUnit_out_ex_exception_3; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_8 = Csr_io_executeUnit_out_ex_exception_8; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_9 = Csr_io_executeUnit_out_ex_exception_9; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_11 = Csr_io_executeUnit_out_ex_exception_11; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_exception_12 = Csr_io_executeUnit_out_ex_exception_12; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_0 = Csr_io_executeUnit_out_ex_interrupt_0; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_1 = Csr_io_executeUnit_out_ex_interrupt_1; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_2 = Csr_io_executeUnit_out_ex_interrupt_2; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_3 = Csr_io_executeUnit_out_ex_interrupt_3; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_4 = Csr_io_executeUnit_out_ex_interrupt_4; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_5 = Csr_io_executeUnit_out_ex_interrupt_5; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_6 = Csr_io_executeUnit_out_ex_interrupt_6; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_7 = Csr_io_executeUnit_out_ex_interrupt_7; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_8 = Csr_io_executeUnit_out_ex_interrupt_8; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_9 = Csr_io_executeUnit_out_ex_interrupt_9; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_10 = Csr_io_executeUnit_out_ex_interrupt_10; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_interrupt_11 = Csr_io_executeUnit_out_ex_interrupt_11; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_tval_1 = Csr_io_executeUnit_out_ex_tval_1; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_tval_2 = Csr_io_executeUnit_out_ex_tval_2; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_ex_tval_12 = Csr_io_executeUnit_out_ex_tval_12; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_flush = Csr_io_executeUnit_out_flush; // @[playground/src/Core.scala 97:19]
  assign ExecuteUnit_io_csr_out_target = Csr_io_executeUnit_out_target; // @[playground/src/Core.scala 97:19]
  assign Csr_clock = clock;
  assign Csr_reset = reset;
  assign Csr_io_ext_int_ei = io_ext_int_ei; // @[playground/src/Core.scala 107:15]
  assign Csr_io_ext_int_ti = io_ext_int_ti; // @[playground/src/Core.scala 107:15]
  assign Csr_io_ext_int_si = io_ext_int_si; // @[playground/src/Core.scala 107:15]
  assign Csr_io_executeUnit_in_valid = ExecuteUnit_io_csr_in_valid; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_pc = ExecuteUnit_io_csr_in_pc; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_info_op = ExecuteUnit_io_csr_in_info_op; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_info_inst = ExecuteUnit_io_csr_in_info_inst; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_src_info_src1_data = ExecuteUnit_io_csr_in_src_info_src1_data; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_1 = ExecuteUnit_io_csr_in_ex_exception_1; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_2 = ExecuteUnit_io_csr_in_ex_exception_2; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_3 = ExecuteUnit_io_csr_in_ex_exception_3; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_8 = ExecuteUnit_io_csr_in_ex_exception_8; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_9 = ExecuteUnit_io_csr_in_ex_exception_9; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_11 = ExecuteUnit_io_csr_in_ex_exception_11; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_exception_12 = ExecuteUnit_io_csr_in_ex_exception_12; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_0 = ExecuteUnit_io_csr_in_ex_interrupt_0; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_1 = ExecuteUnit_io_csr_in_ex_interrupt_1; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_2 = ExecuteUnit_io_csr_in_ex_interrupt_2; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_3 = ExecuteUnit_io_csr_in_ex_interrupt_3; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_4 = ExecuteUnit_io_csr_in_ex_interrupt_4; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_5 = ExecuteUnit_io_csr_in_ex_interrupt_5; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_6 = ExecuteUnit_io_csr_in_ex_interrupt_6; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_7 = ExecuteUnit_io_csr_in_ex_interrupt_7; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_8 = ExecuteUnit_io_csr_in_ex_interrupt_8; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_9 = ExecuteUnit_io_csr_in_ex_interrupt_9; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_10 = ExecuteUnit_io_csr_in_ex_interrupt_10; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_interrupt_11 = ExecuteUnit_io_csr_in_ex_interrupt_11; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_tval_1 = ExecuteUnit_io_csr_in_ex_tval_1; // @[playground/src/Core.scala 97:19]
  assign Csr_io_executeUnit_in_ex_tval_12 = ExecuteUnit_io_csr_in_ex_tval_12; // @[playground/src/Core.scala 97:19]
  assign Csr_io_memoryUnit_in_pc = MemoryUnit_io_csr_in_pc; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_0 = MemoryUnit_io_csr_in_ex_exception_0; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_1 = MemoryUnit_io_csr_in_ex_exception_1; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_2 = MemoryUnit_io_csr_in_ex_exception_2; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_3 = MemoryUnit_io_csr_in_ex_exception_3; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_4 = MemoryUnit_io_csr_in_ex_exception_4; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_5 = MemoryUnit_io_csr_in_ex_exception_5; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_6 = MemoryUnit_io_csr_in_ex_exception_6; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_7 = MemoryUnit_io_csr_in_ex_exception_7; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_8 = MemoryUnit_io_csr_in_ex_exception_8; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_9 = MemoryUnit_io_csr_in_ex_exception_9; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_10 = MemoryUnit_io_csr_in_ex_exception_10; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_11 = MemoryUnit_io_csr_in_ex_exception_11; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_12 = MemoryUnit_io_csr_in_ex_exception_12; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_13 = MemoryUnit_io_csr_in_ex_exception_13; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_14 = MemoryUnit_io_csr_in_ex_exception_14; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_exception_15 = MemoryUnit_io_csr_in_ex_exception_15; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_0 = MemoryUnit_io_csr_in_ex_interrupt_0; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_1 = MemoryUnit_io_csr_in_ex_interrupt_1; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_2 = MemoryUnit_io_csr_in_ex_interrupt_2; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_3 = MemoryUnit_io_csr_in_ex_interrupt_3; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_4 = MemoryUnit_io_csr_in_ex_interrupt_4; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_5 = MemoryUnit_io_csr_in_ex_interrupt_5; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_6 = MemoryUnit_io_csr_in_ex_interrupt_6; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_7 = MemoryUnit_io_csr_in_ex_interrupt_7; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_8 = MemoryUnit_io_csr_in_ex_interrupt_8; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_9 = MemoryUnit_io_csr_in_ex_interrupt_9; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_10 = MemoryUnit_io_csr_in_ex_interrupt_10; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_interrupt_11 = MemoryUnit_io_csr_in_ex_interrupt_11; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_0 = MemoryUnit_io_csr_in_ex_tval_0; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_1 = MemoryUnit_io_csr_in_ex_tval_1; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_2 = MemoryUnit_io_csr_in_ex_tval_2; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_3 = MemoryUnit_io_csr_in_ex_tval_3; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_4 = MemoryUnit_io_csr_in_ex_tval_4; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_5 = MemoryUnit_io_csr_in_ex_tval_5; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_6 = MemoryUnit_io_csr_in_ex_tval_6; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_7 = MemoryUnit_io_csr_in_ex_tval_7; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_8 = MemoryUnit_io_csr_in_ex_tval_8; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_9 = MemoryUnit_io_csr_in_ex_tval_9; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_10 = MemoryUnit_io_csr_in_ex_tval_10; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_11 = MemoryUnit_io_csr_in_ex_tval_11; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_12 = MemoryUnit_io_csr_in_ex_tval_12; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_13 = MemoryUnit_io_csr_in_ex_tval_13; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_14 = MemoryUnit_io_csr_in_ex_tval_14; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_ex_tval_15 = MemoryUnit_io_csr_in_ex_tval_15; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_info_valid = MemoryUnit_io_csr_in_info_valid; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_info_fusel = MemoryUnit_io_csr_in_info_fusel; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_info_op = MemoryUnit_io_csr_in_info_op; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_lr_wen = MemoryUnit_io_csr_in_lr_wen; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_lr_wbit = MemoryUnit_io_csr_in_lr_wbit; // @[playground/src/Core.scala 104:18]
  assign Csr_io_memoryUnit_in_lr_waddr = MemoryUnit_io_csr_in_lr_waddr; // @[playground/src/Core.scala 104:18]
  assign MemoryStage_clock = clock;
  assign MemoryStage_reset = reset;
  assign MemoryStage_io_ctrl_allow_to_go = Ctrl_io_memoryUnit_allow_to_go; // @[playground/src/Core.scala 100:32]
  assign MemoryStage_io_ctrl_clear = Ctrl_io_memoryUnit_do_flush; // @[playground/src/Core.scala 101:32]
  assign MemoryStage_io_executeUnit_inst_0_pc = ExecuteUnit_io_memoryStage_inst_0_pc; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_valid = ExecuteUnit_io_memoryStage_inst_0_info_valid; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_fusel = ExecuteUnit_io_memoryStage_inst_0_info_fusel; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_op = ExecuteUnit_io_memoryStage_inst_0_info_op; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_reg_wen = ExecuteUnit_io_memoryStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_reg_waddr = ExecuteUnit_io_memoryStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_imm = ExecuteUnit_io_memoryStage_inst_0_info_imm; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_info_inst = ExecuteUnit_io_memoryStage_inst_0_info_inst; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_rd_info_wdata_0 = ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_rd_info_wdata_2 = ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_rd_info_wdata_3 = ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_rd_info_wdata_5 = ExecuteUnit_io_memoryStage_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_src_info_src1_data = ExecuteUnit_io_memoryStage_inst_0_src_info_src1_data; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_src_info_src2_data = ExecuteUnit_io_memoryStage_inst_0_src_info_src2_data; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_0 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_1 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_2 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_3 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_8 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_9 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_11 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_exception_12 = ExecuteUnit_io_memoryStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_0 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_1 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_2 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_3 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_4 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_5 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_6 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_7 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_8 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_9 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_10 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_interrupt_11 = ExecuteUnit_io_memoryStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_tval_0 = ExecuteUnit_io_memoryStage_inst_0_ex_tval_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_tval_1 = ExecuteUnit_io_memoryStage_inst_0_ex_tval_1; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_tval_2 = ExecuteUnit_io_memoryStage_inst_0_ex_tval_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_0_ex_tval_12 = ExecuteUnit_io_memoryStage_inst_0_ex_tval_12; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_pc = ExecuteUnit_io_memoryStage_inst_1_pc; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_valid = ExecuteUnit_io_memoryStage_inst_1_info_valid; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_fusel = ExecuteUnit_io_memoryStage_inst_1_info_fusel; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_op = ExecuteUnit_io_memoryStage_inst_1_info_op; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_reg_wen = ExecuteUnit_io_memoryStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_reg_waddr = ExecuteUnit_io_memoryStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_imm = ExecuteUnit_io_memoryStage_inst_1_info_imm; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_info_inst = ExecuteUnit_io_memoryStage_inst_1_info_inst; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_rd_info_wdata_0 = ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_rd_info_wdata_2 = ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_rd_info_wdata_3 = ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_rd_info_wdata_5 = ExecuteUnit_io_memoryStage_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_src_info_src1_data = ExecuteUnit_io_memoryStage_inst_1_src_info_src1_data; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_src_info_src2_data = ExecuteUnit_io_memoryStage_inst_1_src_info_src2_data; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_0 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_1 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_2 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_3 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_8 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_9 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_11 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_exception_12 = ExecuteUnit_io_memoryStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_0 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_1 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_2 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_3 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_4 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_5 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_6 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_7 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_8 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_9 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_10 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_interrupt_11 = ExecuteUnit_io_memoryStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_tval_0 = ExecuteUnit_io_memoryStage_inst_1_ex_tval_0; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_tval_1 = ExecuteUnit_io_memoryStage_inst_1_ex_tval_1; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_tval_2 = ExecuteUnit_io_memoryStage_inst_1_ex_tval_2; // @[playground/src/Core.scala 98:27]
  assign MemoryStage_io_executeUnit_inst_1_ex_tval_12 = ExecuteUnit_io_memoryStage_inst_1_ex_tval_12; // @[playground/src/Core.scala 98:27]
  assign MemoryUnit_clock = clock;
  assign MemoryUnit_reset = reset;
  assign MemoryUnit_io_ctrl_allow_to_go = Ctrl_io_memoryUnit_allow_to_go; // @[playground/src/Core.scala 47:19]
  assign MemoryUnit_io_memoryStage_inst_0_pc = MemoryStage_io_memoryUnit_inst_0_pc; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_valid = MemoryStage_io_memoryUnit_inst_0_info_valid; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_fusel = MemoryStage_io_memoryUnit_inst_0_info_fusel; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_op = MemoryStage_io_memoryUnit_inst_0_info_op; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_reg_wen = MemoryStage_io_memoryUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_reg_waddr = MemoryStage_io_memoryUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_imm = MemoryStage_io_memoryUnit_inst_0_info_imm; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_info_inst = MemoryStage_io_memoryUnit_inst_0_info_inst; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_0 = MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_2 = MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_3 = MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_rd_info_wdata_5 = MemoryStage_io_memoryUnit_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_src_info_src1_data = MemoryStage_io_memoryUnit_inst_0_src_info_src1_data; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_src_info_src2_data = MemoryStage_io_memoryUnit_inst_0_src_info_src2_data; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_0 = MemoryStage_io_memoryUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_1 = MemoryStage_io_memoryUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_2 = MemoryStage_io_memoryUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_3 = MemoryStage_io_memoryUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_8 = MemoryStage_io_memoryUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_9 = MemoryStage_io_memoryUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_11 = MemoryStage_io_memoryUnit_inst_0_ex_exception_11; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_exception_12 = MemoryStage_io_memoryUnit_inst_0_ex_exception_12; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_0 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_1 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_2 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_3 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_4 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_5 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_6 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_7 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_8 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_9 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_10 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_interrupt_11 = MemoryStage_io_memoryUnit_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_tval_0 = MemoryStage_io_memoryUnit_inst_0_ex_tval_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_tval_1 = MemoryStage_io_memoryUnit_inst_0_ex_tval_1; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_tval_2 = MemoryStage_io_memoryUnit_inst_0_ex_tval_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_0_ex_tval_12 = MemoryStage_io_memoryUnit_inst_0_ex_tval_12; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_pc = MemoryStage_io_memoryUnit_inst_1_pc; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_valid = MemoryStage_io_memoryUnit_inst_1_info_valid; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_fusel = MemoryStage_io_memoryUnit_inst_1_info_fusel; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_op = MemoryStage_io_memoryUnit_inst_1_info_op; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_reg_wen = MemoryStage_io_memoryUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_reg_waddr = MemoryStage_io_memoryUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_imm = MemoryStage_io_memoryUnit_inst_1_info_imm; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_info_inst = MemoryStage_io_memoryUnit_inst_1_info_inst; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_0 = MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_2 = MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_3 = MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_rd_info_wdata_5 = MemoryStage_io_memoryUnit_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_src_info_src1_data = MemoryStage_io_memoryUnit_inst_1_src_info_src1_data; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_src_info_src2_data = MemoryStage_io_memoryUnit_inst_1_src_info_src2_data; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_0 = MemoryStage_io_memoryUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_1 = MemoryStage_io_memoryUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_2 = MemoryStage_io_memoryUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_3 = MemoryStage_io_memoryUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_8 = MemoryStage_io_memoryUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_9 = MemoryStage_io_memoryUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_11 = MemoryStage_io_memoryUnit_inst_1_ex_exception_11; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_exception_12 = MemoryStage_io_memoryUnit_inst_1_ex_exception_12; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_0 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_1 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_2 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_3 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_4 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_5 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_6 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_7 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_8 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_9 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_10 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_interrupt_11 = MemoryStage_io_memoryUnit_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_tval_0 = MemoryStage_io_memoryUnit_inst_1_ex_tval_0; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_tval_1 = MemoryStage_io_memoryUnit_inst_1_ex_tval_1; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_tval_2 = MemoryStage_io_memoryUnit_inst_1_ex_tval_2; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_memoryStage_inst_1_ex_tval_12 = MemoryStage_io_memoryUnit_inst_1_ex_tval_12; // @[playground/src/Core.scala 103:26]
  assign MemoryUnit_io_csr_out_flush = Csr_io_memoryUnit_out_flush; // @[playground/src/Core.scala 104:18]
  assign MemoryUnit_io_csr_out_target = Csr_io_memoryUnit_out_target; // @[playground/src/Core.scala 104:18]
  assign MemoryUnit_io_csr_out_lr = Csr_io_memoryUnit_out_lr; // @[playground/src/Core.scala 104:18]
  assign MemoryUnit_io_csr_out_lr_addr = Csr_io_memoryUnit_out_lr_addr; // @[playground/src/Core.scala 104:18]
  assign MemoryUnit_io_dataMemory_in_access_fault = io_data_access_fault; // @[playground/src/Core.scala 110:41]
  assign MemoryUnit_io_dataMemory_in_page_fault = io_data_page_fault; // @[playground/src/Core.scala 111:41]
  assign MemoryUnit_io_dataMemory_in_ready = io_data_dcache_ready; // @[playground/src/Core.scala 112:41]
  assign MemoryUnit_io_dataMemory_in_rdata = io_data_rdata; // @[playground/src/Core.scala 109:41]
  assign WriteBackStage_clock = clock;
  assign WriteBackStage_reset = reset;
  assign WriteBackStage_io_ctrl_allow_to_go = Ctrl_io_writeBackUnit_allow_to_go; // @[playground/src/Core.scala 122:35]
  assign WriteBackStage_io_memoryUnit_inst_0_pc = MemoryUnit_io_writeBackStage_inst_0_pc; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_info_valid = MemoryUnit_io_writeBackStage_inst_0_info_valid; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_info_fusel = MemoryUnit_io_writeBackStage_inst_0_info_fusel; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_info_reg_wen = MemoryUnit_io_writeBackStage_inst_0_info_reg_wen; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_info_reg_waddr = MemoryUnit_io_writeBackStage_inst_0_info_reg_waddr; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_0 = MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_0; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_1 = MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_1; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_2 = MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_2; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_3 = MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_3; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_rd_info_wdata_5 = MemoryUnit_io_writeBackStage_inst_0_rd_info_wdata_5; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_0 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_0; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_1 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_1; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_2 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_2; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_3 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_3; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_4 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_4; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_5 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_5; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_6 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_6; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_7 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_7; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_8 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_8; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_9 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_9; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_11 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_11; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_12 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_12; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_13 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_13; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_exception_15 = MemoryUnit_io_writeBackStage_inst_0_ex_exception_15; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_0 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_1 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_2 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_3 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_4 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_5 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_6 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_7 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_8 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_9 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_10 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_10; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_0_ex_interrupt_11 = MemoryUnit_io_writeBackStage_inst_0_ex_interrupt_11; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_pc = MemoryUnit_io_writeBackStage_inst_1_pc; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_info_valid = MemoryUnit_io_writeBackStage_inst_1_info_valid; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_info_fusel = MemoryUnit_io_writeBackStage_inst_1_info_fusel; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_info_reg_wen = MemoryUnit_io_writeBackStage_inst_1_info_reg_wen; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_info_reg_waddr = MemoryUnit_io_writeBackStage_inst_1_info_reg_waddr; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_0 = MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_0; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_1 = MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_1; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_2 = MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_2; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_3 = MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_3; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_rd_info_wdata_5 = MemoryUnit_io_writeBackStage_inst_1_rd_info_wdata_5; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_0 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_0; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_1 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_1; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_2 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_2; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_3 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_3; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_4 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_4; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_5 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_5; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_6 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_6; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_7 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_7; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_8 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_8; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_9 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_9; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_11 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_11; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_12 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_12; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_13 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_13; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_exception_15 = MemoryUnit_io_writeBackStage_inst_1_ex_exception_15; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_0 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_1 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_2 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_3 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_4 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_5 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_6 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_7 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_8 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_9 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_10 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_10; // @[playground/src/Core.scala 121:29]
  assign WriteBackStage_io_memoryUnit_inst_1_ex_interrupt_11 = MemoryUnit_io_writeBackStage_inst_1_ex_interrupt_11; // @[playground/src/Core.scala 121:29]
  assign WriteBackUnit_clock = clock;
  assign WriteBackUnit_io_ctrl_allow_to_go = Ctrl_io_writeBackUnit_allow_to_go; // @[playground/src/Core.scala 126:22]
  assign WriteBackUnit_io_writeBackStage_inst_0_pc = WriteBackStage_io_writeBackUnit_inst_0_pc; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_info_valid = WriteBackStage_io_writeBackUnit_inst_0_info_valid; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_info_fusel = WriteBackStage_io_writeBackUnit_inst_0_info_fusel; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_info_reg_wen = WriteBackStage_io_writeBackUnit_inst_0_info_reg_wen; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_info_reg_waddr = WriteBackStage_io_writeBackUnit_inst_0_info_reg_waddr; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_0 = WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_0
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_1 = WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_1
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_2 = WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_2
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_3 = WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_3
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_rd_info_wdata_5 = WriteBackStage_io_writeBackUnit_inst_0_rd_info_wdata_5
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_0 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_0; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_1 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_1; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_2 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_2; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_3 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_3; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_4 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_4; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_5 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_5; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_6 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_6; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_7 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_7; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_8 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_8; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_9 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_9; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_11 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_11
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_12 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_12
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_13 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_13
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_exception_15 = WriteBackStage_io_writeBackUnit_inst_0_ex_exception_15
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_0 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_0; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_1 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_1; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_2 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_2; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_3 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_3; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_4 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_4; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_5 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_5; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_6 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_6; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_7 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_7; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_8 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_8; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_9 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_9; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_10 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_10
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_0_ex_interrupt_11 = WriteBackStage_io_writeBackUnit_inst_0_ex_interrupt_11
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_pc = WriteBackStage_io_writeBackUnit_inst_1_pc; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_info_valid = WriteBackStage_io_writeBackUnit_inst_1_info_valid; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_info_fusel = WriteBackStage_io_writeBackUnit_inst_1_info_fusel; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_info_reg_wen = WriteBackStage_io_writeBackUnit_inst_1_info_reg_wen; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_info_reg_waddr = WriteBackStage_io_writeBackUnit_inst_1_info_reg_waddr; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_0 = WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_0
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_1 = WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_1
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_2 = WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_2
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_3 = WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_3
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_rd_info_wdata_5 = WriteBackStage_io_writeBackUnit_inst_1_rd_info_wdata_5
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_0 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_0; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_1 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_1; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_2 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_2; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_3 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_3; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_4 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_4; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_5 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_5; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_6 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_6; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_7 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_7; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_8 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_8; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_9 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_9; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_11 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_11
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_12 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_12
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_13 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_13
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_exception_15 = WriteBackStage_io_writeBackUnit_inst_1_ex_exception_15
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_0 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_0; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_1 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_1; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_2 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_2; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_3 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_3; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_4 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_4; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_5 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_5; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_6 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_6; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_7 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_7; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_8 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_8; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_9 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_9; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_10 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_10
    ; // @[playground/src/Core.scala 125:32]
  assign WriteBackUnit_io_writeBackStage_inst_1_ex_interrupt_11 = WriteBackStage_io_writeBackUnit_inst_1_ex_interrupt_11
    ; // @[playground/src/Core.scala 125:32]
  assign Tlb_clock = clock;
  assign Tlb_reset = reset;
  assign Tlb_io_icache_en = io_inst_tlb_en; // @[playground/src/Core.scala 40:14]
  assign Tlb_io_icache_vaddr = io_inst_tlb_vaddr; // @[playground/src/Core.scala 40:14]
  assign Tlb_io_icache_complete_single_request = io_inst_tlb_complete_single_request; // @[playground/src/Core.scala 40:14]
  assign Tlb_io_dcache_en = io_data_tlb_en; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_vaddr = io_data_tlb_vaddr; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_complete_single_request = io_data_tlb_complete_single_request; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_access_type = io_data_tlb_access_type; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_vpn_ready = io_data_tlb_ptw_vpn_ready; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_valid = io_data_tlb_ptw_pte_valid; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_page_fault = io_data_tlb_ptw_pte_bits_page_fault; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_ppn = io_data_tlb_ptw_pte_bits_entry_ppn; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_d = io_data_tlb_ptw_pte_bits_entry_flag_d; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_g = io_data_tlb_ptw_pte_bits_entry_flag_g; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_u = io_data_tlb_ptw_pte_bits_entry_flag_u; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_x = io_data_tlb_ptw_pte_bits_entry_flag_x; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_w = io_data_tlb_ptw_pte_bits_entry_flag_w; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_r = io_data_tlb_ptw_pte_bits_entry_flag_r; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_entry_flag_v = io_data_tlb_ptw_pte_bits_entry_flag_v; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_dcache_ptw_pte_bits_rmask = io_data_tlb_ptw_pte_bits_rmask; // @[playground/src/Core.scala 41:14]
  assign Tlb_io_csr_satp = Csr_io_tlb_satp; // @[playground/src/Core.scala 42:11]
  assign Tlb_io_csr_mstatus = Csr_io_tlb_mstatus; // @[playground/src/Core.scala 42:11]
  assign Tlb_io_csr_imode = Csr_io_tlb_imode; // @[playground/src/Core.scala 42:11]
  assign Tlb_io_csr_dmode = Csr_io_tlb_dmode; // @[playground/src/Core.scala 42:11]
  assign Tlb_io_sfence_vma_valid = MemoryUnit_io_ctrl_sfence_vma_valid; // @[playground/src/Core.scala 43:18]
  assign Tlb_io_sfence_vma_src_info_src1_data = MemoryUnit_io_ctrl_sfence_vma_src_info_src1_data; // @[playground/src/Core.scala 43:18]
  assign Tlb_io_sfence_vma_src_info_src2_data = MemoryUnit_io_ctrl_sfence_vma_src_info_src2_data; // @[playground/src/Core.scala 43:18]
endmodule
module SimpleDualPortRam(
  input         clock,
  input         reset,
  input  [5:0]  io_raddr, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  output [63:0] io_rdata, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input  [5:0]  io_waddr, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input         io_wen, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input         io_wstrb, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input  [63:0] io_wdata // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] bank [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire  bank_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire [5:0] bank_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire [63:0] bank_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire [63:0] bank_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire [5:0] bank_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire  bank_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  wire  bank_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  reg  bank_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[playground/src/cache/memory/SimpleDualPortRam.scala 69:20]
  assign bank_io_rdata_MPORT_en = bank_io_rdata_MPORT_en_pipe_0;
  assign bank_io_rdata_MPORT_addr = bank_io_rdata_MPORT_addr_pipe_0;
  assign bank_io_rdata_MPORT_data = bank[bank_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
  assign bank_MPORT_data = io_wdata;
  assign bank_MPORT_addr = io_waddr;
  assign bank_MPORT_mask = 1'h1;
  assign bank_MPORT_en = io_wen;
  assign io_rdata = bank_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 85:20 86:18 88:18]
  always @(posedge clock) begin
    if (bank_MPORT_en & bank_MPORT_mask) begin
      bank[bank_MPORT_addr] <= bank_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 83:29]
    end
    bank_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:68 assert(\n"
            ); // @[playground/src/cache/memory/SimpleDualPortRam.scala 68:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fatal; // @[playground/src/cache/memory/SimpleDualPortRam.scala 68:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_io_rdata_MPORT_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LUTRam(
  input         clock,
  input         reset,
  input  [5:0]  io_raddr, // @[playground/src/cache/memory/LUTRam.scala 18:14]
  output [19:0] io_rdata, // @[playground/src/cache/memory/LUTRam.scala 18:14]
  input  [5:0]  io_waddr, // @[playground/src/cache/memory/LUTRam.scala 18:14]
  input  [19:0] io_wdata, // @[playground/src/cache/memory/LUTRam.scala 18:14]
  input         io_wen // @[playground/src/cache/memory/LUTRam.scala 18:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] bank_0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_1; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_2; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_3; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_4; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_5; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_6; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_7; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_8; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_9; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_10; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_11; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_12; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_13; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_14; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_15; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_16; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_17; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_18; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_19; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_20; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_21; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_22; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_23; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_24; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_25; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_26; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_27; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_28; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_29; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_30; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_31; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_32; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_33; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_34; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_35; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_36; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_37; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_38; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_39; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_40; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_41; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_42; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_43; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_44; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_45; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_46; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_47; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_48; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_49; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_50; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_51; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_52; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_53; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_54; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_55; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_56; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_57; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_58; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_59; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_60; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_61; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_62; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  reg [19:0] bank_63; // @[playground/src/cache/memory/LUTRam.scala 55:23]
  wire [19:0] _GEN_1 = 6'h1 == io_raddr ? bank_1 : bank_0; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_2 = 6'h2 == io_raddr ? bank_2 : _GEN_1; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_3 = 6'h3 == io_raddr ? bank_3 : _GEN_2; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_4 = 6'h4 == io_raddr ? bank_4 : _GEN_3; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_5 = 6'h5 == io_raddr ? bank_5 : _GEN_4; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_6 = 6'h6 == io_raddr ? bank_6 : _GEN_5; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_7 = 6'h7 == io_raddr ? bank_7 : _GEN_6; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_8 = 6'h8 == io_raddr ? bank_8 : _GEN_7; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_9 = 6'h9 == io_raddr ? bank_9 : _GEN_8; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_10 = 6'ha == io_raddr ? bank_10 : _GEN_9; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_11 = 6'hb == io_raddr ? bank_11 : _GEN_10; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_12 = 6'hc == io_raddr ? bank_12 : _GEN_11; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_13 = 6'hd == io_raddr ? bank_13 : _GEN_12; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_14 = 6'he == io_raddr ? bank_14 : _GEN_13; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_15 = 6'hf == io_raddr ? bank_15 : _GEN_14; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_16 = 6'h10 == io_raddr ? bank_16 : _GEN_15; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_17 = 6'h11 == io_raddr ? bank_17 : _GEN_16; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_18 = 6'h12 == io_raddr ? bank_18 : _GEN_17; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_19 = 6'h13 == io_raddr ? bank_19 : _GEN_18; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_20 = 6'h14 == io_raddr ? bank_20 : _GEN_19; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_21 = 6'h15 == io_raddr ? bank_21 : _GEN_20; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_22 = 6'h16 == io_raddr ? bank_22 : _GEN_21; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_23 = 6'h17 == io_raddr ? bank_23 : _GEN_22; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_24 = 6'h18 == io_raddr ? bank_24 : _GEN_23; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_25 = 6'h19 == io_raddr ? bank_25 : _GEN_24; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_26 = 6'h1a == io_raddr ? bank_26 : _GEN_25; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_27 = 6'h1b == io_raddr ? bank_27 : _GEN_26; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_28 = 6'h1c == io_raddr ? bank_28 : _GEN_27; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_29 = 6'h1d == io_raddr ? bank_29 : _GEN_28; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_30 = 6'h1e == io_raddr ? bank_30 : _GEN_29; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_31 = 6'h1f == io_raddr ? bank_31 : _GEN_30; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_32 = 6'h20 == io_raddr ? bank_32 : _GEN_31; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_33 = 6'h21 == io_raddr ? bank_33 : _GEN_32; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_34 = 6'h22 == io_raddr ? bank_34 : _GEN_33; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_35 = 6'h23 == io_raddr ? bank_35 : _GEN_34; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_36 = 6'h24 == io_raddr ? bank_36 : _GEN_35; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_37 = 6'h25 == io_raddr ? bank_37 : _GEN_36; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_38 = 6'h26 == io_raddr ? bank_38 : _GEN_37; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_39 = 6'h27 == io_raddr ? bank_39 : _GEN_38; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_40 = 6'h28 == io_raddr ? bank_40 : _GEN_39; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_41 = 6'h29 == io_raddr ? bank_41 : _GEN_40; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_42 = 6'h2a == io_raddr ? bank_42 : _GEN_41; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_43 = 6'h2b == io_raddr ? bank_43 : _GEN_42; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_44 = 6'h2c == io_raddr ? bank_44 : _GEN_43; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_45 = 6'h2d == io_raddr ? bank_45 : _GEN_44; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_46 = 6'h2e == io_raddr ? bank_46 : _GEN_45; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_47 = 6'h2f == io_raddr ? bank_47 : _GEN_46; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_48 = 6'h30 == io_raddr ? bank_48 : _GEN_47; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_49 = 6'h31 == io_raddr ? bank_49 : _GEN_48; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_50 = 6'h32 == io_raddr ? bank_50 : _GEN_49; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_51 = 6'h33 == io_raddr ? bank_51 : _GEN_50; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_52 = 6'h34 == io_raddr ? bank_52 : _GEN_51; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_53 = 6'h35 == io_raddr ? bank_53 : _GEN_52; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_54 = 6'h36 == io_raddr ? bank_54 : _GEN_53; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_55 = 6'h37 == io_raddr ? bank_55 : _GEN_54; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_56 = 6'h38 == io_raddr ? bank_56 : _GEN_55; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_57 = 6'h39 == io_raddr ? bank_57 : _GEN_56; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_58 = 6'h3a == io_raddr ? bank_58 : _GEN_57; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_59 = 6'h3b == io_raddr ? bank_59 : _GEN_58; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_60 = 6'h3c == io_raddr ? bank_60 : _GEN_59; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_61 = 6'h3d == io_raddr ? bank_61 : _GEN_60; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  wire [19:0] _GEN_62 = 6'h3e == io_raddr ? bank_62 : _GEN_61; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  assign io_rdata = 6'h3f == io_raddr ? bank_63 : _GEN_62; // @[playground/src/cache/memory/LUTRam.scala 56:{20,20}]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_0 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h0 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_0 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_1 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_1 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_2 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_2 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_3 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_3 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_4 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h4 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_4 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_5 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h5 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_5 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_6 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h6 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_6 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_7 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h7 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_7 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_8 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h8 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_8 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_9 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h9 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_9 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_10 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'ha == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_10 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_11 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'hb == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_11 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_12 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'hc == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_12 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_13 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'hd == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_13 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_14 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'he == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_14 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_15 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'hf == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_15 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_16 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h10 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_16 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_17 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h11 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_17 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_18 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h12 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_18 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_19 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h13 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_19 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_20 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h14 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_20 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_21 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h15 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_21 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_22 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h16 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_22 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_23 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h17 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_23 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_24 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h18 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_24 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_25 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h19 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_25 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_26 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1a == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_26 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_27 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1b == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_27 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_28 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1c == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_28 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_29 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1d == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_29 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_30 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1e == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_30 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_31 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h1f == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_31 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_32 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h20 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_32 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_33 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h21 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_33 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_34 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h22 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_34 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_35 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h23 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_35 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_36 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h24 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_36 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_37 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h25 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_37 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_38 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h26 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_38 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_39 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h27 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_39 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_40 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h28 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_40 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_41 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h29 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_41 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_42 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2a == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_42 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_43 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2b == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_43 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_44 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2c == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_44 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_45 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2d == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_45 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_46 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2e == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_46 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_47 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h2f == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_47 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_48 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h30 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_48 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_49 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h31 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_49 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_50 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h32 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_50 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_51 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h33 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_51 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_52 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h34 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_52 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_53 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h35 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_53 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_54 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h36 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_54 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_55 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h37 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_55 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_56 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h38 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_56 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_57 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h39 == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_57 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_58 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3a == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_58 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_59 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3b == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_59 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_60 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3c == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_60 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_61 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3d == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_61 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_62 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3e == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_62 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
    if (reset) begin // @[playground/src/cache/memory/LUTRam.scala 55:23]
      bank_63 <= 20'h0; // @[playground/src/cache/memory/LUTRam.scala 55:23]
    end else if (io_wen) begin // @[playground/src/cache/memory/LUTRam.scala 58:18]
      if (6'h3f == io_waddr) begin // @[playground/src/cache/memory/LUTRam.scala 59:22]
        bank_63 <= io_wdata; // @[playground/src/cache/memory/LUTRam.scala 59:22]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bank_0 = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  bank_1 = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  bank_2 = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  bank_3 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  bank_4 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  bank_5 = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  bank_6 = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  bank_7 = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  bank_8 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  bank_9 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  bank_10 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  bank_11 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  bank_12 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  bank_13 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  bank_14 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  bank_15 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  bank_16 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  bank_17 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  bank_18 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  bank_19 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  bank_20 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  bank_21 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  bank_22 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  bank_23 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  bank_24 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  bank_25 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  bank_26 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  bank_27 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  bank_28 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  bank_29 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  bank_30 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  bank_31 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  bank_32 = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  bank_33 = _RAND_33[19:0];
  _RAND_34 = {1{`RANDOM}};
  bank_34 = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  bank_35 = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  bank_36 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  bank_37 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  bank_38 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  bank_39 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  bank_40 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  bank_41 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  bank_42 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  bank_43 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  bank_44 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  bank_45 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  bank_46 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  bank_47 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  bank_48 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  bank_49 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  bank_50 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  bank_51 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  bank_52 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  bank_53 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  bank_54 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  bank_55 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  bank_56 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  bank_57 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  bank_58 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  bank_59 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  bank_60 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  bank_61 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  bank_62 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  bank_63 = _RAND_63[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input         clock,
  input         reset,
  input         io_cpu_req, // @[playground/src/cache/ICache.scala 72:14]
  input         io_cpu_complete_single_request, // @[playground/src/cache/ICache.scala 72:14]
  input  [63:0] io_cpu_addr_0, // @[playground/src/cache/ICache.scala 72:14]
  input  [63:0] io_cpu_addr_1, // @[playground/src/cache/ICache.scala 72:14]
  input         io_cpu_fence_i, // @[playground/src/cache/ICache.scala 72:14]
  input         io_cpu_dcache_stall, // @[playground/src/cache/ICache.scala 72:14]
  output [63:0] io_cpu_inst_0, // @[playground/src/cache/ICache.scala 72:14]
  output [63:0] io_cpu_inst_1, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_inst_valid_0, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_inst_valid_1, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_access_fault, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_page_fault, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_addr_misaligned, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_icache_stall, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_tlb_en, // @[playground/src/cache/ICache.scala 72:14]
  output [63:0] io_cpu_tlb_vaddr, // @[playground/src/cache/ICache.scala 72:14]
  output        io_cpu_tlb_complete_single_request, // @[playground/src/cache/ICache.scala 72:14]
  input         io_cpu_tlb_uncached, // @[playground/src/cache/ICache.scala 72:14]
  input         io_cpu_tlb_hit, // @[playground/src/cache/ICache.scala 72:14]
  input  [19:0] io_cpu_tlb_ptag, // @[playground/src/cache/ICache.scala 72:14]
  input  [31:0] io_cpu_tlb_paddr, // @[playground/src/cache/ICache.scala 72:14]
  input         io_cpu_tlb_page_fault, // @[playground/src/cache/ICache.scala 72:14]
  input         io_axi_ar_ready, // @[playground/src/cache/ICache.scala 72:14]
  output        io_axi_ar_valid, // @[playground/src/cache/ICache.scala 72:14]
  output [31:0] io_axi_ar_bits_addr, // @[playground/src/cache/ICache.scala 72:14]
  output [7:0]  io_axi_ar_bits_len, // @[playground/src/cache/ICache.scala 72:14]
  output [2:0]  io_axi_ar_bits_size, // @[playground/src/cache/ICache.scala 72:14]
  output        io_axi_r_ready, // @[playground/src/cache/ICache.scala 72:14]
  input         io_axi_r_valid, // @[playground/src/cache/ICache.scala 72:14]
  input  [63:0] io_axi_r_bits_data, // @[playground/src/cache/ICache.scala 72:14]
  input  [1:0]  io_axi_r_bits_resp, // @[playground/src/cache/ICache.scala 72:14]
  input         io_axi_r_bits_last // @[playground/src/cache/ICache.scala 72:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
`endif // RANDOMIZE_REG_INIT
  wire  bank_0_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_0_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_0_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_0_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_0_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_1_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_1_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_1_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_1_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_2_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_2_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_2_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_2_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_3_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_3_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_3_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_3_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_4_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_4_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_4_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_4_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_5_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_5_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_5_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_5_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_6_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_6_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_6_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_6_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_7_0_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_7_0_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_7_0_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_7_0_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_0_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_0_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_0_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_0_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_0_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_1_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_1_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_1_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_1_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_1_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_2_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_2_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_2_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_2_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_2_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_3_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_3_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_3_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_3_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_3_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_4_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_4_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_4_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_4_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_4_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_5_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_5_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_5_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_5_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_5_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_6_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_6_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_6_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_6_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_6_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_1_clock; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_1_reset; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_7_0_1_io_raddr; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_7_0_1_io_rdata; // @[playground/src/cache/ICache.scala 168:17]
  wire [5:0] bank_7_0_1_io_waddr; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_1_io_wen; // @[playground/src/cache/ICache.scala 168:17]
  wire  bank_7_0_1_io_wstrb; // @[playground/src/cache/ICache.scala 168:17]
  wire [63:0] bank_7_0_1_io_wdata; // @[playground/src/cache/ICache.scala 168:17]
  wire  tagBram_clock; // @[playground/src/cache/ICache.scala 192:25]
  wire  tagBram_reset; // @[playground/src/cache/ICache.scala 192:25]
  wire [5:0] tagBram_io_raddr; // @[playground/src/cache/ICache.scala 192:25]
  wire [19:0] tagBram_io_rdata; // @[playground/src/cache/ICache.scala 192:25]
  wire [5:0] tagBram_io_waddr; // @[playground/src/cache/ICache.scala 192:25]
  wire [19:0] tagBram_io_wdata; // @[playground/src/cache/ICache.scala 192:25]
  wire  tagBram_io_wen; // @[playground/src/cache/ICache.scala 192:25]
  wire  tagBram_1_clock; // @[playground/src/cache/ICache.scala 192:25]
  wire  tagBram_1_reset; // @[playground/src/cache/ICache.scala 192:25]
  wire [5:0] tagBram_1_io_raddr; // @[playground/src/cache/ICache.scala 192:25]
  wire [19:0] tagBram_1_io_rdata; // @[playground/src/cache/ICache.scala 192:25]
  wire [5:0] tagBram_1_io_waddr; // @[playground/src/cache/ICache.scala 192:25]
  wire [19:0] tagBram_1_io_wdata; // @[playground/src/cache/ICache.scala 192:25]
  wire  tagBram_1_io_wen; // @[playground/src/cache/ICache.scala 192:25]
  wire [2:0] bank_index = io_cpu_addr_0[5:3]; // @[playground/src/cache/ICache.scala 87:35]
  wire  bank_offset = io_cpu_addr_0[2]; // @[playground/src/cache/ICache.scala 88:35]
  reg [2:0] state; // @[playground/src/cache/ICache.scala 92:94]
  reg  valid_0_0; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_1; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_2; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_3; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_4; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_5; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_6; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_7; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_8; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_9; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_10; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_11; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_12; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_13; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_14; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_15; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_16; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_17; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_18; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_19; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_20; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_21; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_22; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_23; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_24; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_25; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_26; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_27; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_28; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_29; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_30; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_31; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_32; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_33; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_34; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_35; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_36; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_37; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_38; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_39; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_40; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_41; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_42; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_43; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_44; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_45; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_46; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_47; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_48; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_49; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_50; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_51; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_52; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_53; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_54; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_55; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_56; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_57; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_58; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_59; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_60; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_61; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_62; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_0_63; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_0; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_1; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_2; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_3; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_4; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_5; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_6; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_7; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_8; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_9; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_10; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_11; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_12; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_13; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_14; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_15; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_16; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_17; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_18; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_19; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_20; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_21; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_22; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_23; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_24; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_25; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_26; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_27; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_28; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_29; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_30; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_31; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_32; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_33; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_34; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_35; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_36; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_37; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_38; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_39; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_40; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_41; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_42; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_43; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_44; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_45; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_46; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_47; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_48; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_49; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_50; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_51; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_52; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_53; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_54; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_55; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_56; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_57; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_58; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_59; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_60; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_61; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_62; // @[playground/src/cache/ICache.scala 95:22]
  reg  valid_1_63; // @[playground/src/cache/ICache.scala 95:22]
  wire  _use_next_addr_T = state == 3'h0; // @[playground/src/cache/ICache.scala 98:30]
  wire  use_next_addr = state == 3'h0 | state == 3'h3; // @[playground/src/cache/ICache.scala 98:42]
  wire [63:0] _GEN_1 = use_next_addr ? io_cpu_addr_1 : io_cpu_addr_0; // @[playground/src/cache/ICache.scala 102:{47,47}]
  reg [19:0] tag_0; // @[playground/src/cache/ICache.scala 104:26]
  reg [19:0] tag_1; // @[playground/src/cache/ICache.scala 104:26]
  reg  tag_wstrb_0; // @[playground/src/cache/ICache.scala 106:26]
  reg  tag_wstrb_1; // @[playground/src/cache/ICache.scala 106:26]
  reg [19:0] tag_wdata; // @[playground/src/cache/ICache.scala 107:26]
  reg  lru_0; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_1; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_2; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_3; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_4; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_5; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_6; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_7; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_8; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_9; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_10; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_11; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_12; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_13; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_14; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_15; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_16; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_17; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_18; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_19; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_20; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_21; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_22; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_23; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_24; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_25; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_26; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_27; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_28; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_29; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_30; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_31; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_32; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_33; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_34; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_35; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_36; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_37; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_38; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_39; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_40; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_41; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_42; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_43; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_44; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_45; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_46; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_47; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_48; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_49; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_50; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_51; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_52; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_53; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_54; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_55; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_56; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_57; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_58; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_59; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_60; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_61; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_62; // @[playground/src/cache/ICache.scala 110:20]
  reg  lru_63; // @[playground/src/cache/ICache.scala 110:20]
  wire [5:0] replace_index = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  reg  replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 117:30]
  reg  replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 117:30]
  wire  _GEN_3 = 6'h1 == replace_index ? valid_0_1 : valid_0_0; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_4 = 6'h2 == replace_index ? valid_0_2 : _GEN_3; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_5 = 6'h3 == replace_index ? valid_0_3 : _GEN_4; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_6 = 6'h4 == replace_index ? valid_0_4 : _GEN_5; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_7 = 6'h5 == replace_index ? valid_0_5 : _GEN_6; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_8 = 6'h6 == replace_index ? valid_0_6 : _GEN_7; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_9 = 6'h7 == replace_index ? valid_0_7 : _GEN_8; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_10 = 6'h8 == replace_index ? valid_0_8 : _GEN_9; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_11 = 6'h9 == replace_index ? valid_0_9 : _GEN_10; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_12 = 6'ha == replace_index ? valid_0_10 : _GEN_11; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_13 = 6'hb == replace_index ? valid_0_11 : _GEN_12; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_14 = 6'hc == replace_index ? valid_0_12 : _GEN_13; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_15 = 6'hd == replace_index ? valid_0_13 : _GEN_14; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_16 = 6'he == replace_index ? valid_0_14 : _GEN_15; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_17 = 6'hf == replace_index ? valid_0_15 : _GEN_16; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_18 = 6'h10 == replace_index ? valid_0_16 : _GEN_17; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_19 = 6'h11 == replace_index ? valid_0_17 : _GEN_18; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_20 = 6'h12 == replace_index ? valid_0_18 : _GEN_19; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_21 = 6'h13 == replace_index ? valid_0_19 : _GEN_20; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_22 = 6'h14 == replace_index ? valid_0_20 : _GEN_21; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_23 = 6'h15 == replace_index ? valid_0_21 : _GEN_22; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_24 = 6'h16 == replace_index ? valid_0_22 : _GEN_23; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_25 = 6'h17 == replace_index ? valid_0_23 : _GEN_24; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_26 = 6'h18 == replace_index ? valid_0_24 : _GEN_25; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_27 = 6'h19 == replace_index ? valid_0_25 : _GEN_26; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_28 = 6'h1a == replace_index ? valid_0_26 : _GEN_27; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_29 = 6'h1b == replace_index ? valid_0_27 : _GEN_28; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_30 = 6'h1c == replace_index ? valid_0_28 : _GEN_29; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_31 = 6'h1d == replace_index ? valid_0_29 : _GEN_30; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_32 = 6'h1e == replace_index ? valid_0_30 : _GEN_31; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_33 = 6'h1f == replace_index ? valid_0_31 : _GEN_32; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_34 = 6'h20 == replace_index ? valid_0_32 : _GEN_33; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_35 = 6'h21 == replace_index ? valid_0_33 : _GEN_34; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_36 = 6'h22 == replace_index ? valid_0_34 : _GEN_35; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_37 = 6'h23 == replace_index ? valid_0_35 : _GEN_36; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_38 = 6'h24 == replace_index ? valid_0_36 : _GEN_37; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_39 = 6'h25 == replace_index ? valid_0_37 : _GEN_38; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_40 = 6'h26 == replace_index ? valid_0_38 : _GEN_39; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_41 = 6'h27 == replace_index ? valid_0_39 : _GEN_40; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_42 = 6'h28 == replace_index ? valid_0_40 : _GEN_41; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_43 = 6'h29 == replace_index ? valid_0_41 : _GEN_42; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_44 = 6'h2a == replace_index ? valid_0_42 : _GEN_43; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_45 = 6'h2b == replace_index ? valid_0_43 : _GEN_44; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_46 = 6'h2c == replace_index ? valid_0_44 : _GEN_45; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_47 = 6'h2d == replace_index ? valid_0_45 : _GEN_46; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_48 = 6'h2e == replace_index ? valid_0_46 : _GEN_47; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_49 = 6'h2f == replace_index ? valid_0_47 : _GEN_48; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_50 = 6'h30 == replace_index ? valid_0_48 : _GEN_49; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_51 = 6'h31 == replace_index ? valid_0_49 : _GEN_50; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_52 = 6'h32 == replace_index ? valid_0_50 : _GEN_51; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_53 = 6'h33 == replace_index ? valid_0_51 : _GEN_52; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_54 = 6'h34 == replace_index ? valid_0_52 : _GEN_53; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_55 = 6'h35 == replace_index ? valid_0_53 : _GEN_54; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_56 = 6'h36 == replace_index ? valid_0_54 : _GEN_55; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_57 = 6'h37 == replace_index ? valid_0_55 : _GEN_56; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_58 = 6'h38 == replace_index ? valid_0_56 : _GEN_57; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_59 = 6'h39 == replace_index ? valid_0_57 : _GEN_58; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_60 = 6'h3a == replace_index ? valid_0_58 : _GEN_59; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_61 = 6'h3b == replace_index ? valid_0_59 : _GEN_60; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_62 = 6'h3c == replace_index ? valid_0_60 : _GEN_61; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_63 = 6'h3d == replace_index ? valid_0_61 : _GEN_62; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_64 = 6'h3e == replace_index ? valid_0_62 : _GEN_63; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_65 = 6'h3f == replace_index ? valid_0_63 : _GEN_64; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  tag_compare_valid_0 = tag_0 == io_cpu_tlb_ptag & _GEN_65; // @[playground/src/cache/ICache.scala 122:88]
  wire  _GEN_67 = 6'h1 == replace_index ? valid_1_1 : valid_1_0; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_68 = 6'h2 == replace_index ? valid_1_2 : _GEN_67; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_69 = 6'h3 == replace_index ? valid_1_3 : _GEN_68; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_70 = 6'h4 == replace_index ? valid_1_4 : _GEN_69; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_71 = 6'h5 == replace_index ? valid_1_5 : _GEN_70; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_72 = 6'h6 == replace_index ? valid_1_6 : _GEN_71; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_73 = 6'h7 == replace_index ? valid_1_7 : _GEN_72; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_74 = 6'h8 == replace_index ? valid_1_8 : _GEN_73; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_75 = 6'h9 == replace_index ? valid_1_9 : _GEN_74; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_76 = 6'ha == replace_index ? valid_1_10 : _GEN_75; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_77 = 6'hb == replace_index ? valid_1_11 : _GEN_76; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_78 = 6'hc == replace_index ? valid_1_12 : _GEN_77; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_79 = 6'hd == replace_index ? valid_1_13 : _GEN_78; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_80 = 6'he == replace_index ? valid_1_14 : _GEN_79; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_81 = 6'hf == replace_index ? valid_1_15 : _GEN_80; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_82 = 6'h10 == replace_index ? valid_1_16 : _GEN_81; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_83 = 6'h11 == replace_index ? valid_1_17 : _GEN_82; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_84 = 6'h12 == replace_index ? valid_1_18 : _GEN_83; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_85 = 6'h13 == replace_index ? valid_1_19 : _GEN_84; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_86 = 6'h14 == replace_index ? valid_1_20 : _GEN_85; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_87 = 6'h15 == replace_index ? valid_1_21 : _GEN_86; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_88 = 6'h16 == replace_index ? valid_1_22 : _GEN_87; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_89 = 6'h17 == replace_index ? valid_1_23 : _GEN_88; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_90 = 6'h18 == replace_index ? valid_1_24 : _GEN_89; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_91 = 6'h19 == replace_index ? valid_1_25 : _GEN_90; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_92 = 6'h1a == replace_index ? valid_1_26 : _GEN_91; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_93 = 6'h1b == replace_index ? valid_1_27 : _GEN_92; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_94 = 6'h1c == replace_index ? valid_1_28 : _GEN_93; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_95 = 6'h1d == replace_index ? valid_1_29 : _GEN_94; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_96 = 6'h1e == replace_index ? valid_1_30 : _GEN_95; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_97 = 6'h1f == replace_index ? valid_1_31 : _GEN_96; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_98 = 6'h20 == replace_index ? valid_1_32 : _GEN_97; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_99 = 6'h21 == replace_index ? valid_1_33 : _GEN_98; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_100 = 6'h22 == replace_index ? valid_1_34 : _GEN_99; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_101 = 6'h23 == replace_index ? valid_1_35 : _GEN_100; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_102 = 6'h24 == replace_index ? valid_1_36 : _GEN_101; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_103 = 6'h25 == replace_index ? valid_1_37 : _GEN_102; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_104 = 6'h26 == replace_index ? valid_1_38 : _GEN_103; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_105 = 6'h27 == replace_index ? valid_1_39 : _GEN_104; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_106 = 6'h28 == replace_index ? valid_1_40 : _GEN_105; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_107 = 6'h29 == replace_index ? valid_1_41 : _GEN_106; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_108 = 6'h2a == replace_index ? valid_1_42 : _GEN_107; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_109 = 6'h2b == replace_index ? valid_1_43 : _GEN_108; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_110 = 6'h2c == replace_index ? valid_1_44 : _GEN_109; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_111 = 6'h2d == replace_index ? valid_1_45 : _GEN_110; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_112 = 6'h2e == replace_index ? valid_1_46 : _GEN_111; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_113 = 6'h2f == replace_index ? valid_1_47 : _GEN_112; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_114 = 6'h30 == replace_index ? valid_1_48 : _GEN_113; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_115 = 6'h31 == replace_index ? valid_1_49 : _GEN_114; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_116 = 6'h32 == replace_index ? valid_1_50 : _GEN_115; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_117 = 6'h33 == replace_index ? valid_1_51 : _GEN_116; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_118 = 6'h34 == replace_index ? valid_1_52 : _GEN_117; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_119 = 6'h35 == replace_index ? valid_1_53 : _GEN_118; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_120 = 6'h36 == replace_index ? valid_1_54 : _GEN_119; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_121 = 6'h37 == replace_index ? valid_1_55 : _GEN_120; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_122 = 6'h38 == replace_index ? valid_1_56 : _GEN_121; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_123 = 6'h39 == replace_index ? valid_1_57 : _GEN_122; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_124 = 6'h3a == replace_index ? valid_1_58 : _GEN_123; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_125 = 6'h3b == replace_index ? valid_1_59 : _GEN_124; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_126 = 6'h3c == replace_index ? valid_1_60 : _GEN_125; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_127 = 6'h3d == replace_index ? valid_1_61 : _GEN_126; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_128 = 6'h3e == replace_index ? valid_1_62 : _GEN_127; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  _GEN_129 = 6'h3f == replace_index ? valid_1_63 : _GEN_128; // @[playground/src/cache/ICache.scala 122:{88,88}]
  wire  tag_compare_valid_1 = tag_1 == io_cpu_tlb_ptag & _GEN_129; // @[playground/src/cache/ICache.scala 122:88]
  wire  cache_hit = tag_compare_valid_0 | tag_compare_valid_1; // @[playground/src/cache/ICache.scala 123:55]
  wire  cache_hit_available = cache_hit & io_cpu_tlb_hit & ~io_cpu_tlb_uncached; // @[playground/src/cache/ICache.scala 124:57]
  wire [63:0] data_0_0_0 = bank_0_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] data_0_1_0 = bank_1_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire  _GEN_2165 = ~tag_compare_valid_1; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] _GEN_131 = ~tag_compare_valid_1 & 3'h1 == bank_index ? data_0_1_0 : data_0_0_0; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_0_2_0 = bank_2_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_132 = ~tag_compare_valid_1 & 3'h2 == bank_index ? data_0_2_0 : _GEN_131; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_0_3_0 = bank_3_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_133 = ~tag_compare_valid_1 & 3'h3 == bank_index ? data_0_3_0 : _GEN_132; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_0_4_0 = bank_4_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_134 = ~tag_compare_valid_1 & 3'h4 == bank_index ? data_0_4_0 : _GEN_133; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_0_5_0 = bank_5_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_135 = ~tag_compare_valid_1 & 3'h5 == bank_index ? data_0_5_0 : _GEN_134; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_0_6_0 = bank_6_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_136 = ~tag_compare_valid_1 & 3'h6 == bank_index ? data_0_6_0 : _GEN_135; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_0_7_0 = bank_7_0_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_137 = ~tag_compare_valid_1 & 3'h7 == bank_index ? data_0_7_0 : _GEN_136; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_0_0 = bank_0_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_138 = tag_compare_valid_1 & 3'h0 == bank_index ? data_1_0_0 : _GEN_137; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_1_0 = bank_1_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_139 = tag_compare_valid_1 & 3'h1 == bank_index ? data_1_1_0 : _GEN_138; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_2_0 = bank_2_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_140 = tag_compare_valid_1 & 3'h2 == bank_index ? data_1_2_0 : _GEN_139; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_3_0 = bank_3_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_141 = tag_compare_valid_1 & 3'h3 == bank_index ? data_1_3_0 : _GEN_140; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_4_0 = bank_4_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_142 = tag_compare_valid_1 & 3'h4 == bank_index ? data_1_4_0 : _GEN_141; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_5_0 = bank_5_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_143 = tag_compare_valid_1 & 3'h5 == bank_index ? data_1_5_0 : _GEN_142; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_6_0 = bank_6_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_144 = tag_compare_valid_1 & 3'h6 == bank_index ? data_1_6_0 : _GEN_143; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [63:0] data_1_7_0 = bank_7_0_1_io_rdata; // @[playground/src/cache/ICache.scala 101:25 175:29]
  wire [63:0] _GEN_145 = tag_compare_valid_1 & 3'h7 == bank_index ? data_1_7_0 : _GEN_144; // @[playground/src/cache/ICache.scala 129:{72,72}]
  wire [31:0] inst_in_bank_0 = _GEN_145[31:0]; // @[playground/src/cache/ICache.scala 129:72]
  wire [31:0] inst_in_bank_1 = _GEN_145[63:32]; // @[playground/src/cache/ICache.scala 129:72]
  wire [1:0] _inst_T_3 = {{1'd0}, bank_offset}; // @[playground/src/cache/ICache.scala 140:26]
  wire [31:0] inst_0 = _inst_T_3[0] ? inst_in_bank_1 : inst_in_bank_0; // @[playground/src/cache/ICache.scala 138:{10,10}]
  wire  _inst_T_8 = 1'h1 <= 1'h1 - bank_offset; // @[playground/src/cache/ICache.scala 139:13]
  wire  _inst_T_10 = 1'h1 + bank_offset; // @[playground/src/cache/ICache.scala 140:26]
  wire [31:0] _GEN_149 = _inst_T_10 ? inst_in_bank_1 : inst_in_bank_0; // @[playground/src/cache/ICache.scala 138:{10,10}]
  wire [31:0] inst_1 = _inst_T_8 ? _GEN_149 : 32'h0; // @[playground/src/cache/ICache.scala 138:10]
  wire  inst_valid_1 = cache_hit_available & _inst_T_8; // @[playground/src/cache/ICache.scala 146:57]
  reg [31:0] rdata_in_wait_0_inst; // @[playground/src/cache/ICache.scala 149:30]
  reg  rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 149:30]
  reg [31:0] rdata_in_wait_1_inst; // @[playground/src/cache/ICache.scala 149:30]
  reg  rdata_in_wait_1_valid; // @[playground/src/cache/ICache.scala 149:30]
  wire  _io_cpu_inst_valid_0_T_1 = _use_next_addr_T ? cache_hit_available : rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 186:32]
  wire [31:0] _io_cpu_inst_0_T_1 = _use_next_addr_T ? inst_0 : rdata_in_wait_0_inst; // @[playground/src/cache/ICache.scala 187:32]
  wire  _io_cpu_inst_valid_1_T_1 = _use_next_addr_T ? inst_valid_1 : rdata_in_wait_1_valid; // @[playground/src/cache/ICache.scala 186:32]
  wire [31:0] _io_cpu_inst_1_T_1 = _use_next_addr_T ? inst_1 : rdata_in_wait_1_inst; // @[playground/src/cache/ICache.scala 187:32]
  reg [31:0] ar_addr; // @[playground/src/cache/ICache.scala 207:24]
  reg [7:0] ar_len; // @[playground/src/cache/ICache.scala 207:24]
  reg [2:0] ar_size; // @[playground/src/cache/ICache.scala 207:24]
  reg  arvalid; // @[playground/src/cache/ICache.scala 208:24]
  reg  rready; // @[playground/src/cache/ICache.scala 213:23]
  reg  access_fault; // @[playground/src/cache/ICache.scala 217:32]
  reg  page_fault; // @[playground/src/cache/ICache.scala 218:32]
  reg  addr_misaligned; // @[playground/src/cache/ICache.scala 219:32]
  wire  _addr_err_T_27 = _GEN_1[39] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_29 = _GEN_1[40] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_31 = _GEN_1[41] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_33 = _GEN_1[42] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_35 = _GEN_1[43] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_37 = _GEN_1[44] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_39 = _GEN_1[45] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_41 = _GEN_1[46] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_43 = _GEN_1[47] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_45 = _GEN_1[48] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_47 = _GEN_1[49] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_49 = _GEN_1[50] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_51 = _GEN_1[51] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_53 = _GEN_1[52] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_55 = _GEN_1[53] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_57 = _GEN_1[54] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_59 = _GEN_1[55] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_61 = _GEN_1[56] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_63 = _GEN_1[57] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_65 = _GEN_1[58] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_67 = _GEN_1[59] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_69 = _GEN_1[60] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_71 = _GEN_1[61] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_73 = _GEN_1[62] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_75 = _GEN_1[63] != _GEN_1[38]; // @[playground/src/cache/ICache.scala 225:14]
  wire  _addr_err_T_101 = |_GEN_1[1:0]; // @[playground/src/cache/ICache.scala 227:65]
  wire  addr_err = _addr_err_T_27 | _addr_err_T_29 | _addr_err_T_31 | _addr_err_T_33 | _addr_err_T_35 | _addr_err_T_37
     | _addr_err_T_39 | _addr_err_T_41 | _addr_err_T_43 | _addr_err_T_45 | _addr_err_T_47 | _addr_err_T_49 |
    _addr_err_T_51 | _addr_err_T_53 | _addr_err_T_55 | _addr_err_T_57 | _addr_err_T_59 | _addr_err_T_61 | _addr_err_T_63
     | _addr_err_T_65 | _addr_err_T_67 | _addr_err_T_69 | _addr_err_T_71 | _addr_err_T_73 | _addr_err_T_75 |
    _addr_err_T_101; // @[playground/src/cache/ICache.scala 226:23]
  wire  _GEN_151 = _addr_err_T_101 ? 1'h0 : 1'h1; // @[playground/src/cache/ICache.scala 235:23 240:79 243:26]
  wire [31:0] _ar_addr_T_1 = {io_cpu_tlb_paddr[31:6],6'h0}; // @[playground/src/cache/ICache.scala 259:25]
  wire  _GEN_153 = 6'h1 == replace_index ? lru_1 : lru_0; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_154 = 6'h2 == replace_index ? lru_2 : _GEN_153; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_155 = 6'h3 == replace_index ? lru_3 : _GEN_154; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_156 = 6'h4 == replace_index ? lru_4 : _GEN_155; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_157 = 6'h5 == replace_index ? lru_5 : _GEN_156; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_158 = 6'h6 == replace_index ? lru_6 : _GEN_157; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_159 = 6'h7 == replace_index ? lru_7 : _GEN_158; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_160 = 6'h8 == replace_index ? lru_8 : _GEN_159; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_161 = 6'h9 == replace_index ? lru_9 : _GEN_160; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_162 = 6'ha == replace_index ? lru_10 : _GEN_161; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_163 = 6'hb == replace_index ? lru_11 : _GEN_162; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_164 = 6'hc == replace_index ? lru_12 : _GEN_163; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_165 = 6'hd == replace_index ? lru_13 : _GEN_164; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_166 = 6'he == replace_index ? lru_14 : _GEN_165; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_167 = 6'hf == replace_index ? lru_15 : _GEN_166; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_168 = 6'h10 == replace_index ? lru_16 : _GEN_167; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_169 = 6'h11 == replace_index ? lru_17 : _GEN_168; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_170 = 6'h12 == replace_index ? lru_18 : _GEN_169; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_171 = 6'h13 == replace_index ? lru_19 : _GEN_170; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_172 = 6'h14 == replace_index ? lru_20 : _GEN_171; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_173 = 6'h15 == replace_index ? lru_21 : _GEN_172; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_174 = 6'h16 == replace_index ? lru_22 : _GEN_173; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_175 = 6'h17 == replace_index ? lru_23 : _GEN_174; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_176 = 6'h18 == replace_index ? lru_24 : _GEN_175; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_177 = 6'h19 == replace_index ? lru_25 : _GEN_176; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_178 = 6'h1a == replace_index ? lru_26 : _GEN_177; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_179 = 6'h1b == replace_index ? lru_27 : _GEN_178; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_180 = 6'h1c == replace_index ? lru_28 : _GEN_179; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_181 = 6'h1d == replace_index ? lru_29 : _GEN_180; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_182 = 6'h1e == replace_index ? lru_30 : _GEN_181; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_183 = 6'h1f == replace_index ? lru_31 : _GEN_182; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_184 = 6'h20 == replace_index ? lru_32 : _GEN_183; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_185 = 6'h21 == replace_index ? lru_33 : _GEN_184; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_186 = 6'h22 == replace_index ? lru_34 : _GEN_185; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_187 = 6'h23 == replace_index ? lru_35 : _GEN_186; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_188 = 6'h24 == replace_index ? lru_36 : _GEN_187; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_189 = 6'h25 == replace_index ? lru_37 : _GEN_188; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_190 = 6'h26 == replace_index ? lru_38 : _GEN_189; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_191 = 6'h27 == replace_index ? lru_39 : _GEN_190; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_192 = 6'h28 == replace_index ? lru_40 : _GEN_191; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_193 = 6'h29 == replace_index ? lru_41 : _GEN_192; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_194 = 6'h2a == replace_index ? lru_42 : _GEN_193; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_195 = 6'h2b == replace_index ? lru_43 : _GEN_194; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_196 = 6'h2c == replace_index ? lru_44 : _GEN_195; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_197 = 6'h2d == replace_index ? lru_45 : _GEN_196; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_198 = 6'h2e == replace_index ? lru_46 : _GEN_197; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_199 = 6'h2f == replace_index ? lru_47 : _GEN_198; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_200 = 6'h30 == replace_index ? lru_48 : _GEN_199; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_201 = 6'h31 == replace_index ? lru_49 : _GEN_200; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_202 = 6'h32 == replace_index ? lru_50 : _GEN_201; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_203 = 6'h33 == replace_index ? lru_51 : _GEN_202; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_204 = 6'h34 == replace_index ? lru_52 : _GEN_203; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_205 = 6'h35 == replace_index ? lru_53 : _GEN_204; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_206 = 6'h36 == replace_index ? lru_54 : _GEN_205; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_207 = 6'h37 == replace_index ? lru_55 : _GEN_206; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_208 = 6'h38 == replace_index ? lru_56 : _GEN_207; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_209 = 6'h39 == replace_index ? lru_57 : _GEN_208; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_210 = 6'h3a == replace_index ? lru_58 : _GEN_209; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_211 = 6'h3b == replace_index ? lru_59 : _GEN_210; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_212 = 6'h3c == replace_index ? lru_60 : _GEN_211; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_213 = 6'h3d == replace_index ? lru_61 : _GEN_212; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_214 = 6'h3e == replace_index ? lru_62 : _GEN_213; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_215 = 6'h3f == replace_index ? lru_63 : _GEN_214; // @[playground/src/cache/ICache.scala 264:{50,50}]
  wire  _GEN_216 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_217 = _GEN_215 ? 1'h0 : replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_218 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_219 = _GEN_215 ? 1'h0 : replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_220 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_221 = _GEN_215 ? 1'h0 : replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_222 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_223 = _GEN_215 ? 1'h0 : replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_224 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_225 = _GEN_215 ? 1'h0 : replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_226 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_227 = _GEN_215 ? 1'h0 : replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_228 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_229 = _GEN_215 ? 1'h0 : replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_230 = ~_GEN_215 ? 1'h0 : replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_231 = _GEN_215 ? 1'h0 : replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 117:30 264:{50,50}]
  wire  _GEN_2187 = ~_GEN_215; // @[playground/src/cache/ICache.scala 265:{45,45}]
  wire  _GEN_232 = ~_GEN_215 | _GEN_216; // @[playground/src/cache/ICache.scala 265:{45,45}]
  wire  _GEN_233 = _GEN_215 | _GEN_217; // @[playground/src/cache/ICache.scala 265:{45,45}]
  wire  _GEN_234 = _GEN_2187 | tag_wstrb_0; // @[playground/src/cache/ICache.scala 106:26 266:{45,45}]
  wire  _GEN_235 = _GEN_215 | tag_wstrb_1; // @[playground/src/cache/ICache.scala 106:26 266:{45,45}]
  wire  _GEN_236 = _GEN_2187 & 6'h0 == replace_index | valid_0_0; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_237 = _GEN_2187 & 6'h1 == replace_index | valid_0_1; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_238 = _GEN_2187 & 6'h2 == replace_index | valid_0_2; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_239 = _GEN_2187 & 6'h3 == replace_index | valid_0_3; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_240 = _GEN_2187 & 6'h4 == replace_index | valid_0_4; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_241 = _GEN_2187 & 6'h5 == replace_index | valid_0_5; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_242 = _GEN_2187 & 6'h6 == replace_index | valid_0_6; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_243 = _GEN_2187 & 6'h7 == replace_index | valid_0_7; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_244 = _GEN_2187 & 6'h8 == replace_index | valid_0_8; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_245 = _GEN_2187 & 6'h9 == replace_index | valid_0_9; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_246 = _GEN_2187 & 6'ha == replace_index | valid_0_10; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_247 = _GEN_2187 & 6'hb == replace_index | valid_0_11; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_248 = _GEN_2187 & 6'hc == replace_index | valid_0_12; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_249 = _GEN_2187 & 6'hd == replace_index | valid_0_13; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_250 = _GEN_2187 & 6'he == replace_index | valid_0_14; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_251 = _GEN_2187 & 6'hf == replace_index | valid_0_15; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_252 = _GEN_2187 & 6'h10 == replace_index | valid_0_16; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_253 = _GEN_2187 & 6'h11 == replace_index | valid_0_17; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_254 = _GEN_2187 & 6'h12 == replace_index | valid_0_18; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_255 = _GEN_2187 & 6'h13 == replace_index | valid_0_19; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_256 = _GEN_2187 & 6'h14 == replace_index | valid_0_20; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_257 = _GEN_2187 & 6'h15 == replace_index | valid_0_21; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_258 = _GEN_2187 & 6'h16 == replace_index | valid_0_22; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_259 = _GEN_2187 & 6'h17 == replace_index | valid_0_23; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_260 = _GEN_2187 & 6'h18 == replace_index | valid_0_24; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_261 = _GEN_2187 & 6'h19 == replace_index | valid_0_25; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_262 = _GEN_2187 & 6'h1a == replace_index | valid_0_26; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_263 = _GEN_2187 & 6'h1b == replace_index | valid_0_27; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_264 = _GEN_2187 & 6'h1c == replace_index | valid_0_28; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_265 = _GEN_2187 & 6'h1d == replace_index | valid_0_29; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_266 = _GEN_2187 & 6'h1e == replace_index | valid_0_30; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_267 = _GEN_2187 & 6'h1f == replace_index | valid_0_31; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_268 = _GEN_2187 & 6'h20 == replace_index | valid_0_32; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_269 = _GEN_2187 & 6'h21 == replace_index | valid_0_33; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_270 = _GEN_2187 & 6'h22 == replace_index | valid_0_34; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_271 = _GEN_2187 & 6'h23 == replace_index | valid_0_35; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_272 = _GEN_2187 & 6'h24 == replace_index | valid_0_36; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_273 = _GEN_2187 & 6'h25 == replace_index | valid_0_37; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_274 = _GEN_2187 & 6'h26 == replace_index | valid_0_38; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_275 = _GEN_2187 & 6'h27 == replace_index | valid_0_39; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_276 = _GEN_2187 & 6'h28 == replace_index | valid_0_40; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_277 = _GEN_2187 & 6'h29 == replace_index | valid_0_41; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_278 = _GEN_2187 & 6'h2a == replace_index | valid_0_42; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_279 = _GEN_2187 & 6'h2b == replace_index | valid_0_43; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_280 = _GEN_2187 & 6'h2c == replace_index | valid_0_44; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_281 = _GEN_2187 & 6'h2d == replace_index | valid_0_45; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_282 = _GEN_2187 & 6'h2e == replace_index | valid_0_46; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_283 = _GEN_2187 & 6'h2f == replace_index | valid_0_47; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_284 = _GEN_2187 & 6'h30 == replace_index | valid_0_48; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_285 = _GEN_2187 & 6'h31 == replace_index | valid_0_49; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_286 = _GEN_2187 & 6'h32 == replace_index | valid_0_50; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_287 = _GEN_2187 & 6'h33 == replace_index | valid_0_51; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_288 = _GEN_2187 & 6'h34 == replace_index | valid_0_52; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_289 = _GEN_2187 & 6'h35 == replace_index | valid_0_53; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_290 = _GEN_2187 & 6'h36 == replace_index | valid_0_54; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_291 = _GEN_2187 & 6'h37 == replace_index | valid_0_55; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_292 = _GEN_2187 & 6'h38 == replace_index | valid_0_56; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_293 = _GEN_2187 & 6'h39 == replace_index | valid_0_57; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_294 = _GEN_2187 & 6'h3a == replace_index | valid_0_58; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_295 = _GEN_2187 & 6'h3b == replace_index | valid_0_59; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_296 = _GEN_2187 & 6'h3c == replace_index | valid_0_60; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_297 = _GEN_2187 & 6'h3d == replace_index | valid_0_61; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_298 = _GEN_2187 & 6'h3e == replace_index | valid_0_62; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_299 = _GEN_2187 & 6'h3f == replace_index | valid_0_63; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_300 = _GEN_215 & 6'h0 == replace_index | valid_1_0; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_301 = _GEN_215 & 6'h1 == replace_index | valid_1_1; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_302 = _GEN_215 & 6'h2 == replace_index | valid_1_2; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_303 = _GEN_215 & 6'h3 == replace_index | valid_1_3; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_304 = _GEN_215 & 6'h4 == replace_index | valid_1_4; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_305 = _GEN_215 & 6'h5 == replace_index | valid_1_5; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_306 = _GEN_215 & 6'h6 == replace_index | valid_1_6; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_307 = _GEN_215 & 6'h7 == replace_index | valid_1_7; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_308 = _GEN_215 & 6'h8 == replace_index | valid_1_8; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_309 = _GEN_215 & 6'h9 == replace_index | valid_1_9; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_310 = _GEN_215 & 6'ha == replace_index | valid_1_10; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_311 = _GEN_215 & 6'hb == replace_index | valid_1_11; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_312 = _GEN_215 & 6'hc == replace_index | valid_1_12; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_313 = _GEN_215 & 6'hd == replace_index | valid_1_13; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_314 = _GEN_215 & 6'he == replace_index | valid_1_14; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_315 = _GEN_215 & 6'hf == replace_index | valid_1_15; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_316 = _GEN_215 & 6'h10 == replace_index | valid_1_16; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_317 = _GEN_215 & 6'h11 == replace_index | valid_1_17; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_318 = _GEN_215 & 6'h12 == replace_index | valid_1_18; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_319 = _GEN_215 & 6'h13 == replace_index | valid_1_19; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_320 = _GEN_215 & 6'h14 == replace_index | valid_1_20; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_321 = _GEN_215 & 6'h15 == replace_index | valid_1_21; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_322 = _GEN_215 & 6'h16 == replace_index | valid_1_22; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_323 = _GEN_215 & 6'h17 == replace_index | valid_1_23; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_324 = _GEN_215 & 6'h18 == replace_index | valid_1_24; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_325 = _GEN_215 & 6'h19 == replace_index | valid_1_25; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_326 = _GEN_215 & 6'h1a == replace_index | valid_1_26; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_327 = _GEN_215 & 6'h1b == replace_index | valid_1_27; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_328 = _GEN_215 & 6'h1c == replace_index | valid_1_28; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_329 = _GEN_215 & 6'h1d == replace_index | valid_1_29; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_330 = _GEN_215 & 6'h1e == replace_index | valid_1_30; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_331 = _GEN_215 & 6'h1f == replace_index | valid_1_31; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_332 = _GEN_215 & 6'h20 == replace_index | valid_1_32; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_333 = _GEN_215 & 6'h21 == replace_index | valid_1_33; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_334 = _GEN_215 & 6'h22 == replace_index | valid_1_34; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_335 = _GEN_215 & 6'h23 == replace_index | valid_1_35; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_336 = _GEN_215 & 6'h24 == replace_index | valid_1_36; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_337 = _GEN_215 & 6'h25 == replace_index | valid_1_37; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_338 = _GEN_215 & 6'h26 == replace_index | valid_1_38; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_339 = _GEN_215 & 6'h27 == replace_index | valid_1_39; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_340 = _GEN_215 & 6'h28 == replace_index | valid_1_40; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_341 = _GEN_215 & 6'h29 == replace_index | valid_1_41; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_342 = _GEN_215 & 6'h2a == replace_index | valid_1_42; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_343 = _GEN_215 & 6'h2b == replace_index | valid_1_43; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_344 = _GEN_215 & 6'h2c == replace_index | valid_1_44; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_345 = _GEN_215 & 6'h2d == replace_index | valid_1_45; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_346 = _GEN_215 & 6'h2e == replace_index | valid_1_46; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_347 = _GEN_215 & 6'h2f == replace_index | valid_1_47; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_348 = _GEN_215 & 6'h30 == replace_index | valid_1_48; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_349 = _GEN_215 & 6'h31 == replace_index | valid_1_49; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_350 = _GEN_215 & 6'h32 == replace_index | valid_1_50; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_351 = _GEN_215 & 6'h33 == replace_index | valid_1_51; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_352 = _GEN_215 & 6'h34 == replace_index | valid_1_52; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_353 = _GEN_215 & 6'h35 == replace_index | valid_1_53; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_354 = _GEN_215 & 6'h36 == replace_index | valid_1_54; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_355 = _GEN_215 & 6'h37 == replace_index | valid_1_55; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_356 = _GEN_215 & 6'h38 == replace_index | valid_1_56; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_357 = _GEN_215 & 6'h39 == replace_index | valid_1_57; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_358 = _GEN_215 & 6'h3a == replace_index | valid_1_58; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_359 = _GEN_215 & 6'h3b == replace_index | valid_1_59; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_360 = _GEN_215 & 6'h3c == replace_index | valid_1_60; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_361 = _GEN_215 & 6'h3d == replace_index | valid_1_61; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_362 = _GEN_215 & 6'h3e == replace_index | valid_1_62; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_363 = _GEN_215 & 6'h3f == replace_index | valid_1_63; // @[playground/src/cache/ICache.scala 268:{45,45} 95:22]
  wire  _GEN_364 = 6'h0 == replace_index ? _GEN_2165 : lru_0; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_365 = 6'h1 == replace_index ? _GEN_2165 : lru_1; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_366 = 6'h2 == replace_index ? _GEN_2165 : lru_2; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_367 = 6'h3 == replace_index ? _GEN_2165 : lru_3; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_368 = 6'h4 == replace_index ? _GEN_2165 : lru_4; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_369 = 6'h5 == replace_index ? _GEN_2165 : lru_5; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_370 = 6'h6 == replace_index ? _GEN_2165 : lru_6; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_371 = 6'h7 == replace_index ? _GEN_2165 : lru_7; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_372 = 6'h8 == replace_index ? _GEN_2165 : lru_8; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_373 = 6'h9 == replace_index ? _GEN_2165 : lru_9; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_374 = 6'ha == replace_index ? _GEN_2165 : lru_10; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_375 = 6'hb == replace_index ? _GEN_2165 : lru_11; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_376 = 6'hc == replace_index ? _GEN_2165 : lru_12; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_377 = 6'hd == replace_index ? _GEN_2165 : lru_13; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_378 = 6'he == replace_index ? _GEN_2165 : lru_14; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_379 = 6'hf == replace_index ? _GEN_2165 : lru_15; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_380 = 6'h10 == replace_index ? _GEN_2165 : lru_16; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_381 = 6'h11 == replace_index ? _GEN_2165 : lru_17; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_382 = 6'h12 == replace_index ? _GEN_2165 : lru_18; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_383 = 6'h13 == replace_index ? _GEN_2165 : lru_19; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_384 = 6'h14 == replace_index ? _GEN_2165 : lru_20; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_385 = 6'h15 == replace_index ? _GEN_2165 : lru_21; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_386 = 6'h16 == replace_index ? _GEN_2165 : lru_22; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_387 = 6'h17 == replace_index ? _GEN_2165 : lru_23; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_388 = 6'h18 == replace_index ? _GEN_2165 : lru_24; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_389 = 6'h19 == replace_index ? _GEN_2165 : lru_25; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_390 = 6'h1a == replace_index ? _GEN_2165 : lru_26; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_391 = 6'h1b == replace_index ? _GEN_2165 : lru_27; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_392 = 6'h1c == replace_index ? _GEN_2165 : lru_28; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_393 = 6'h1d == replace_index ? _GEN_2165 : lru_29; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_394 = 6'h1e == replace_index ? _GEN_2165 : lru_30; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_395 = 6'h1f == replace_index ? _GEN_2165 : lru_31; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_396 = 6'h20 == replace_index ? _GEN_2165 : lru_32; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_397 = 6'h21 == replace_index ? _GEN_2165 : lru_33; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_398 = 6'h22 == replace_index ? _GEN_2165 : lru_34; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_399 = 6'h23 == replace_index ? _GEN_2165 : lru_35; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_400 = 6'h24 == replace_index ? _GEN_2165 : lru_36; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_401 = 6'h25 == replace_index ? _GEN_2165 : lru_37; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_402 = 6'h26 == replace_index ? _GEN_2165 : lru_38; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_403 = 6'h27 == replace_index ? _GEN_2165 : lru_39; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_404 = 6'h28 == replace_index ? _GEN_2165 : lru_40; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_405 = 6'h29 == replace_index ? _GEN_2165 : lru_41; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_406 = 6'h2a == replace_index ? _GEN_2165 : lru_42; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_407 = 6'h2b == replace_index ? _GEN_2165 : lru_43; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_408 = 6'h2c == replace_index ? _GEN_2165 : lru_44; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_409 = 6'h2d == replace_index ? _GEN_2165 : lru_45; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_410 = 6'h2e == replace_index ? _GEN_2165 : lru_46; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_411 = 6'h2f == replace_index ? _GEN_2165 : lru_47; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_412 = 6'h30 == replace_index ? _GEN_2165 : lru_48; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_413 = 6'h31 == replace_index ? _GEN_2165 : lru_49; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_414 = 6'h32 == replace_index ? _GEN_2165 : lru_50; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_415 = 6'h33 == replace_index ? _GEN_2165 : lru_51; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_416 = 6'h34 == replace_index ? _GEN_2165 : lru_52; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_417 = 6'h35 == replace_index ? _GEN_2165 : lru_53; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_418 = 6'h36 == replace_index ? _GEN_2165 : lru_54; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_419 = 6'h37 == replace_index ? _GEN_2165 : lru_55; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_420 = 6'h38 == replace_index ? _GEN_2165 : lru_56; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_421 = 6'h39 == replace_index ? _GEN_2165 : lru_57; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_422 = 6'h3a == replace_index ? _GEN_2165 : lru_58; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_423 = 6'h3b == replace_index ? _GEN_2165 : lru_59; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_424 = 6'h3c == replace_index ? _GEN_2165 : lru_60; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_425 = 6'h3d == replace_index ? _GEN_2165 : lru_61; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_426 = 6'h3e == replace_index ? _GEN_2165 : lru_62; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire  _GEN_427 = 6'h3f == replace_index ? _GEN_2165 : lru_63; // @[playground/src/cache/ICache.scala 110:20 270:{23,23}]
  wire [2:0] _GEN_428 = ~io_cpu_complete_single_request ? 3'h3 : state; // @[playground/src/cache/ICache.scala 271:49 272:19 92:94]
  wire [31:0] _GEN_429 = ~io_cpu_complete_single_request ? inst_1 : rdata_in_wait_1_inst; // @[playground/src/cache/ICache.scala 149:30 271:49 273:71]
  wire  _GEN_430 = ~io_cpu_complete_single_request ? cache_hit_available : rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 149:30 271:49 274:72]
  wire  _GEN_431 = ~io_cpu_complete_single_request ? inst_valid_1 : rdata_in_wait_1_valid; // @[playground/src/cache/ICache.scala 149:30 271:49 274:72]
  wire  _GEN_432 = ~io_cpu_icache_stall ? _GEN_364 : lru_0; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_433 = ~io_cpu_icache_stall ? _GEN_365 : lru_1; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_434 = ~io_cpu_icache_stall ? _GEN_366 : lru_2; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_435 = ~io_cpu_icache_stall ? _GEN_367 : lru_3; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_436 = ~io_cpu_icache_stall ? _GEN_368 : lru_4; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_437 = ~io_cpu_icache_stall ? _GEN_369 : lru_5; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_438 = ~io_cpu_icache_stall ? _GEN_370 : lru_6; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_439 = ~io_cpu_icache_stall ? _GEN_371 : lru_7; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_440 = ~io_cpu_icache_stall ? _GEN_372 : lru_8; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_441 = ~io_cpu_icache_stall ? _GEN_373 : lru_9; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_442 = ~io_cpu_icache_stall ? _GEN_374 : lru_10; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_443 = ~io_cpu_icache_stall ? _GEN_375 : lru_11; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_444 = ~io_cpu_icache_stall ? _GEN_376 : lru_12; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_445 = ~io_cpu_icache_stall ? _GEN_377 : lru_13; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_446 = ~io_cpu_icache_stall ? _GEN_378 : lru_14; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_447 = ~io_cpu_icache_stall ? _GEN_379 : lru_15; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_448 = ~io_cpu_icache_stall ? _GEN_380 : lru_16; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_449 = ~io_cpu_icache_stall ? _GEN_381 : lru_17; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_450 = ~io_cpu_icache_stall ? _GEN_382 : lru_18; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_451 = ~io_cpu_icache_stall ? _GEN_383 : lru_19; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_452 = ~io_cpu_icache_stall ? _GEN_384 : lru_20; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_453 = ~io_cpu_icache_stall ? _GEN_385 : lru_21; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_454 = ~io_cpu_icache_stall ? _GEN_386 : lru_22; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_455 = ~io_cpu_icache_stall ? _GEN_387 : lru_23; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_456 = ~io_cpu_icache_stall ? _GEN_388 : lru_24; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_457 = ~io_cpu_icache_stall ? _GEN_389 : lru_25; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_458 = ~io_cpu_icache_stall ? _GEN_390 : lru_26; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_459 = ~io_cpu_icache_stall ? _GEN_391 : lru_27; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_460 = ~io_cpu_icache_stall ? _GEN_392 : lru_28; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_461 = ~io_cpu_icache_stall ? _GEN_393 : lru_29; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_462 = ~io_cpu_icache_stall ? _GEN_394 : lru_30; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_463 = ~io_cpu_icache_stall ? _GEN_395 : lru_31; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_464 = ~io_cpu_icache_stall ? _GEN_396 : lru_32; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_465 = ~io_cpu_icache_stall ? _GEN_397 : lru_33; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_466 = ~io_cpu_icache_stall ? _GEN_398 : lru_34; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_467 = ~io_cpu_icache_stall ? _GEN_399 : lru_35; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_468 = ~io_cpu_icache_stall ? _GEN_400 : lru_36; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_469 = ~io_cpu_icache_stall ? _GEN_401 : lru_37; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_470 = ~io_cpu_icache_stall ? _GEN_402 : lru_38; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_471 = ~io_cpu_icache_stall ? _GEN_403 : lru_39; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_472 = ~io_cpu_icache_stall ? _GEN_404 : lru_40; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_473 = ~io_cpu_icache_stall ? _GEN_405 : lru_41; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_474 = ~io_cpu_icache_stall ? _GEN_406 : lru_42; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_475 = ~io_cpu_icache_stall ? _GEN_407 : lru_43; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_476 = ~io_cpu_icache_stall ? _GEN_408 : lru_44; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_477 = ~io_cpu_icache_stall ? _GEN_409 : lru_45; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_478 = ~io_cpu_icache_stall ? _GEN_410 : lru_46; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_479 = ~io_cpu_icache_stall ? _GEN_411 : lru_47; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_480 = ~io_cpu_icache_stall ? _GEN_412 : lru_48; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_481 = ~io_cpu_icache_stall ? _GEN_413 : lru_49; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_482 = ~io_cpu_icache_stall ? _GEN_414 : lru_50; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_483 = ~io_cpu_icache_stall ? _GEN_415 : lru_51; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_484 = ~io_cpu_icache_stall ? _GEN_416 : lru_52; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_485 = ~io_cpu_icache_stall ? _GEN_417 : lru_53; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_486 = ~io_cpu_icache_stall ? _GEN_418 : lru_54; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_487 = ~io_cpu_icache_stall ? _GEN_419 : lru_55; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_488 = ~io_cpu_icache_stall ? _GEN_420 : lru_56; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_489 = ~io_cpu_icache_stall ? _GEN_421 : lru_57; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_490 = ~io_cpu_icache_stall ? _GEN_422 : lru_58; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_491 = ~io_cpu_icache_stall ? _GEN_423 : lru_59; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_492 = ~io_cpu_icache_stall ? _GEN_424 : lru_60; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_493 = ~io_cpu_icache_stall ? _GEN_425 : lru_61; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_494 = ~io_cpu_icache_stall ? _GEN_426 : lru_62; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire  _GEN_495 = ~io_cpu_icache_stall ? _GEN_427 : lru_63; // @[playground/src/cache/ICache.scala 110:20 269:42]
  wire [2:0] _GEN_496 = ~io_cpu_icache_stall ? _GEN_428 : state; // @[playground/src/cache/ICache.scala 269:42 92:94]
  wire [31:0] _GEN_497 = ~io_cpu_icache_stall ? _GEN_429 : rdata_in_wait_1_inst; // @[playground/src/cache/ICache.scala 149:30 269:42]
  wire  _GEN_498 = ~io_cpu_icache_stall ? _GEN_430 : rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 149:30 269:42]
  wire  _GEN_499 = ~io_cpu_icache_stall ? _GEN_431 : rdata_in_wait_1_valid; // @[playground/src/cache/ICache.scala 149:30 269:42]
  wire [2:0] _GEN_500 = ~cache_hit ? 3'h2 : _GEN_496; // @[playground/src/cache/ICache.scala 256:32 257:17]
  wire [31:0] _GEN_501 = ~cache_hit ? _ar_addr_T_1 : ar_addr; // @[playground/src/cache/ICache.scala 256:32 259:19 207:24]
  wire [7:0] _GEN_502 = ~cache_hit ? 8'h7 : ar_len; // @[playground/src/cache/ICache.scala 256:32 260:19 207:24]
  wire [2:0] _GEN_503 = ~cache_hit ? 3'h3 : ar_size; // @[playground/src/cache/ICache.scala 256:32 261:19 207:24]
  wire  _GEN_504 = ~cache_hit | arvalid; // @[playground/src/cache/ICache.scala 256:32 262:19 208:24]
  wire  _GEN_505 = ~cache_hit ? _GEN_232 : replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_506 = ~cache_hit ? _GEN_233 : replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_507 = ~cache_hit ? _GEN_218 : replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_508 = ~cache_hit ? _GEN_219 : replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_509 = ~cache_hit ? _GEN_220 : replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_510 = ~cache_hit ? _GEN_221 : replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_511 = ~cache_hit ? _GEN_222 : replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_512 = ~cache_hit ? _GEN_223 : replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_513 = ~cache_hit ? _GEN_224 : replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_514 = ~cache_hit ? _GEN_225 : replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_515 = ~cache_hit ? _GEN_226 : replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_516 = ~cache_hit ? _GEN_227 : replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_517 = ~cache_hit ? _GEN_228 : replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_518 = ~cache_hit ? _GEN_229 : replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_519 = ~cache_hit ? _GEN_230 : replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_520 = ~cache_hit ? _GEN_231 : replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 117:30 256:32]
  wire  _GEN_521 = ~cache_hit ? _GEN_234 : tag_wstrb_0; // @[playground/src/cache/ICache.scala 106:26 256:32]
  wire  _GEN_522 = ~cache_hit ? _GEN_235 : tag_wstrb_1; // @[playground/src/cache/ICache.scala 106:26 256:32]
  wire [19:0] _GEN_523 = ~cache_hit ? io_cpu_tlb_ptag : tag_wdata; // @[playground/src/cache/ICache.scala 107:26 256:32 267:45]
  wire  _GEN_524 = ~cache_hit ? _GEN_236 : valid_0_0; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_525 = ~cache_hit ? _GEN_237 : valid_0_1; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_526 = ~cache_hit ? _GEN_238 : valid_0_2; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_527 = ~cache_hit ? _GEN_239 : valid_0_3; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_528 = ~cache_hit ? _GEN_240 : valid_0_4; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_529 = ~cache_hit ? _GEN_241 : valid_0_5; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_530 = ~cache_hit ? _GEN_242 : valid_0_6; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_531 = ~cache_hit ? _GEN_243 : valid_0_7; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_532 = ~cache_hit ? _GEN_244 : valid_0_8; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_533 = ~cache_hit ? _GEN_245 : valid_0_9; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_534 = ~cache_hit ? _GEN_246 : valid_0_10; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_535 = ~cache_hit ? _GEN_247 : valid_0_11; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_536 = ~cache_hit ? _GEN_248 : valid_0_12; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_537 = ~cache_hit ? _GEN_249 : valid_0_13; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_538 = ~cache_hit ? _GEN_250 : valid_0_14; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_539 = ~cache_hit ? _GEN_251 : valid_0_15; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_540 = ~cache_hit ? _GEN_252 : valid_0_16; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_541 = ~cache_hit ? _GEN_253 : valid_0_17; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_542 = ~cache_hit ? _GEN_254 : valid_0_18; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_543 = ~cache_hit ? _GEN_255 : valid_0_19; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_544 = ~cache_hit ? _GEN_256 : valid_0_20; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_545 = ~cache_hit ? _GEN_257 : valid_0_21; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_546 = ~cache_hit ? _GEN_258 : valid_0_22; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_547 = ~cache_hit ? _GEN_259 : valid_0_23; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_548 = ~cache_hit ? _GEN_260 : valid_0_24; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_549 = ~cache_hit ? _GEN_261 : valid_0_25; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_550 = ~cache_hit ? _GEN_262 : valid_0_26; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_551 = ~cache_hit ? _GEN_263 : valid_0_27; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_552 = ~cache_hit ? _GEN_264 : valid_0_28; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_553 = ~cache_hit ? _GEN_265 : valid_0_29; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_554 = ~cache_hit ? _GEN_266 : valid_0_30; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_555 = ~cache_hit ? _GEN_267 : valid_0_31; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_556 = ~cache_hit ? _GEN_268 : valid_0_32; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_557 = ~cache_hit ? _GEN_269 : valid_0_33; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_558 = ~cache_hit ? _GEN_270 : valid_0_34; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_559 = ~cache_hit ? _GEN_271 : valid_0_35; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_560 = ~cache_hit ? _GEN_272 : valid_0_36; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_561 = ~cache_hit ? _GEN_273 : valid_0_37; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_562 = ~cache_hit ? _GEN_274 : valid_0_38; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_563 = ~cache_hit ? _GEN_275 : valid_0_39; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_564 = ~cache_hit ? _GEN_276 : valid_0_40; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_565 = ~cache_hit ? _GEN_277 : valid_0_41; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_566 = ~cache_hit ? _GEN_278 : valid_0_42; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_567 = ~cache_hit ? _GEN_279 : valid_0_43; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_568 = ~cache_hit ? _GEN_280 : valid_0_44; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_569 = ~cache_hit ? _GEN_281 : valid_0_45; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_570 = ~cache_hit ? _GEN_282 : valid_0_46; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_571 = ~cache_hit ? _GEN_283 : valid_0_47; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_572 = ~cache_hit ? _GEN_284 : valid_0_48; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_573 = ~cache_hit ? _GEN_285 : valid_0_49; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_574 = ~cache_hit ? _GEN_286 : valid_0_50; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_575 = ~cache_hit ? _GEN_287 : valid_0_51; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_576 = ~cache_hit ? _GEN_288 : valid_0_52; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_577 = ~cache_hit ? _GEN_289 : valid_0_53; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_578 = ~cache_hit ? _GEN_290 : valid_0_54; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_579 = ~cache_hit ? _GEN_291 : valid_0_55; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_580 = ~cache_hit ? _GEN_292 : valid_0_56; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_581 = ~cache_hit ? _GEN_293 : valid_0_57; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_582 = ~cache_hit ? _GEN_294 : valid_0_58; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_583 = ~cache_hit ? _GEN_295 : valid_0_59; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_584 = ~cache_hit ? _GEN_296 : valid_0_60; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_585 = ~cache_hit ? _GEN_297 : valid_0_61; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_586 = ~cache_hit ? _GEN_298 : valid_0_62; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_587 = ~cache_hit ? _GEN_299 : valid_0_63; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_588 = ~cache_hit ? _GEN_300 : valid_1_0; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_589 = ~cache_hit ? _GEN_301 : valid_1_1; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_590 = ~cache_hit ? _GEN_302 : valid_1_2; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_591 = ~cache_hit ? _GEN_303 : valid_1_3; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_592 = ~cache_hit ? _GEN_304 : valid_1_4; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_593 = ~cache_hit ? _GEN_305 : valid_1_5; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_594 = ~cache_hit ? _GEN_306 : valid_1_6; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_595 = ~cache_hit ? _GEN_307 : valid_1_7; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_596 = ~cache_hit ? _GEN_308 : valid_1_8; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_597 = ~cache_hit ? _GEN_309 : valid_1_9; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_598 = ~cache_hit ? _GEN_310 : valid_1_10; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_599 = ~cache_hit ? _GEN_311 : valid_1_11; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_600 = ~cache_hit ? _GEN_312 : valid_1_12; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_601 = ~cache_hit ? _GEN_313 : valid_1_13; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_602 = ~cache_hit ? _GEN_314 : valid_1_14; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_603 = ~cache_hit ? _GEN_315 : valid_1_15; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_604 = ~cache_hit ? _GEN_316 : valid_1_16; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_605 = ~cache_hit ? _GEN_317 : valid_1_17; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_606 = ~cache_hit ? _GEN_318 : valid_1_18; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_607 = ~cache_hit ? _GEN_319 : valid_1_19; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_608 = ~cache_hit ? _GEN_320 : valid_1_20; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_609 = ~cache_hit ? _GEN_321 : valid_1_21; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_610 = ~cache_hit ? _GEN_322 : valid_1_22; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_611 = ~cache_hit ? _GEN_323 : valid_1_23; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_612 = ~cache_hit ? _GEN_324 : valid_1_24; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_613 = ~cache_hit ? _GEN_325 : valid_1_25; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_614 = ~cache_hit ? _GEN_326 : valid_1_26; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_615 = ~cache_hit ? _GEN_327 : valid_1_27; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_616 = ~cache_hit ? _GEN_328 : valid_1_28; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_617 = ~cache_hit ? _GEN_329 : valid_1_29; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_618 = ~cache_hit ? _GEN_330 : valid_1_30; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_619 = ~cache_hit ? _GEN_331 : valid_1_31; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_620 = ~cache_hit ? _GEN_332 : valid_1_32; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_621 = ~cache_hit ? _GEN_333 : valid_1_33; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_622 = ~cache_hit ? _GEN_334 : valid_1_34; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_623 = ~cache_hit ? _GEN_335 : valid_1_35; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_624 = ~cache_hit ? _GEN_336 : valid_1_36; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_625 = ~cache_hit ? _GEN_337 : valid_1_37; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_626 = ~cache_hit ? _GEN_338 : valid_1_38; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_627 = ~cache_hit ? _GEN_339 : valid_1_39; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_628 = ~cache_hit ? _GEN_340 : valid_1_40; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_629 = ~cache_hit ? _GEN_341 : valid_1_41; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_630 = ~cache_hit ? _GEN_342 : valid_1_42; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_631 = ~cache_hit ? _GEN_343 : valid_1_43; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_632 = ~cache_hit ? _GEN_344 : valid_1_44; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_633 = ~cache_hit ? _GEN_345 : valid_1_45; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_634 = ~cache_hit ? _GEN_346 : valid_1_46; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_635 = ~cache_hit ? _GEN_347 : valid_1_47; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_636 = ~cache_hit ? _GEN_348 : valid_1_48; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_637 = ~cache_hit ? _GEN_349 : valid_1_49; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_638 = ~cache_hit ? _GEN_350 : valid_1_50; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_639 = ~cache_hit ? _GEN_351 : valid_1_51; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_640 = ~cache_hit ? _GEN_352 : valid_1_52; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_641 = ~cache_hit ? _GEN_353 : valid_1_53; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_642 = ~cache_hit ? _GEN_354 : valid_1_54; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_643 = ~cache_hit ? _GEN_355 : valid_1_55; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_644 = ~cache_hit ? _GEN_356 : valid_1_56; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_645 = ~cache_hit ? _GEN_357 : valid_1_57; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_646 = ~cache_hit ? _GEN_358 : valid_1_58; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_647 = ~cache_hit ? _GEN_359 : valid_1_59; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_648 = ~cache_hit ? _GEN_360 : valid_1_60; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_649 = ~cache_hit ? _GEN_361 : valid_1_61; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_650 = ~cache_hit ? _GEN_362 : valid_1_62; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_651 = ~cache_hit ? _GEN_363 : valid_1_63; // @[playground/src/cache/ICache.scala 256:32 95:22]
  wire  _GEN_652 = ~cache_hit ? lru_0 : _GEN_432; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_653 = ~cache_hit ? lru_1 : _GEN_433; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_654 = ~cache_hit ? lru_2 : _GEN_434; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_655 = ~cache_hit ? lru_3 : _GEN_435; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_656 = ~cache_hit ? lru_4 : _GEN_436; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_657 = ~cache_hit ? lru_5 : _GEN_437; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_658 = ~cache_hit ? lru_6 : _GEN_438; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_659 = ~cache_hit ? lru_7 : _GEN_439; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_660 = ~cache_hit ? lru_8 : _GEN_440; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_661 = ~cache_hit ? lru_9 : _GEN_441; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_662 = ~cache_hit ? lru_10 : _GEN_442; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_663 = ~cache_hit ? lru_11 : _GEN_443; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_664 = ~cache_hit ? lru_12 : _GEN_444; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_665 = ~cache_hit ? lru_13 : _GEN_445; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_666 = ~cache_hit ? lru_14 : _GEN_446; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_667 = ~cache_hit ? lru_15 : _GEN_447; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_668 = ~cache_hit ? lru_16 : _GEN_448; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_669 = ~cache_hit ? lru_17 : _GEN_449; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_670 = ~cache_hit ? lru_18 : _GEN_450; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_671 = ~cache_hit ? lru_19 : _GEN_451; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_672 = ~cache_hit ? lru_20 : _GEN_452; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_673 = ~cache_hit ? lru_21 : _GEN_453; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_674 = ~cache_hit ? lru_22 : _GEN_454; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_675 = ~cache_hit ? lru_23 : _GEN_455; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_676 = ~cache_hit ? lru_24 : _GEN_456; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_677 = ~cache_hit ? lru_25 : _GEN_457; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_678 = ~cache_hit ? lru_26 : _GEN_458; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_679 = ~cache_hit ? lru_27 : _GEN_459; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_680 = ~cache_hit ? lru_28 : _GEN_460; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_681 = ~cache_hit ? lru_29 : _GEN_461; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_682 = ~cache_hit ? lru_30 : _GEN_462; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_683 = ~cache_hit ? lru_31 : _GEN_463; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_684 = ~cache_hit ? lru_32 : _GEN_464; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_685 = ~cache_hit ? lru_33 : _GEN_465; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_686 = ~cache_hit ? lru_34 : _GEN_466; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_687 = ~cache_hit ? lru_35 : _GEN_467; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_688 = ~cache_hit ? lru_36 : _GEN_468; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_689 = ~cache_hit ? lru_37 : _GEN_469; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_690 = ~cache_hit ? lru_38 : _GEN_470; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_691 = ~cache_hit ? lru_39 : _GEN_471; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_692 = ~cache_hit ? lru_40 : _GEN_472; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_693 = ~cache_hit ? lru_41 : _GEN_473; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_694 = ~cache_hit ? lru_42 : _GEN_474; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_695 = ~cache_hit ? lru_43 : _GEN_475; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_696 = ~cache_hit ? lru_44 : _GEN_476; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_697 = ~cache_hit ? lru_45 : _GEN_477; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_698 = ~cache_hit ? lru_46 : _GEN_478; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_699 = ~cache_hit ? lru_47 : _GEN_479; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_700 = ~cache_hit ? lru_48 : _GEN_480; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_701 = ~cache_hit ? lru_49 : _GEN_481; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_702 = ~cache_hit ? lru_50 : _GEN_482; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_703 = ~cache_hit ? lru_51 : _GEN_483; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_704 = ~cache_hit ? lru_52 : _GEN_484; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_705 = ~cache_hit ? lru_53 : _GEN_485; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_706 = ~cache_hit ? lru_54 : _GEN_486; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_707 = ~cache_hit ? lru_55 : _GEN_487; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_708 = ~cache_hit ? lru_56 : _GEN_488; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_709 = ~cache_hit ? lru_57 : _GEN_489; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_710 = ~cache_hit ? lru_58 : _GEN_490; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_711 = ~cache_hit ? lru_59 : _GEN_491; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_712 = ~cache_hit ? lru_60 : _GEN_492; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_713 = ~cache_hit ? lru_61 : _GEN_493; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_714 = ~cache_hit ? lru_62 : _GEN_494; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire  _GEN_715 = ~cache_hit ? lru_63 : _GEN_495; // @[playground/src/cache/ICache.scala 110:20 256:32]
  wire [31:0] _GEN_716 = ~cache_hit ? rdata_in_wait_1_inst : _GEN_497; // @[playground/src/cache/ICache.scala 149:30 256:32]
  wire  _GEN_717 = ~cache_hit ? rdata_in_wait_0_valid : _GEN_498; // @[playground/src/cache/ICache.scala 149:30 256:32]
  wire  _GEN_718 = ~cache_hit ? rdata_in_wait_1_valid : _GEN_499; // @[playground/src/cache/ICache.scala 149:30 256:32]
  wire [2:0] _GEN_719 = io_cpu_tlb_uncached ? 3'h1 : _GEN_500; // @[playground/src/cache/ICache.scala 250:41 251:19]
  wire [31:0] _GEN_720 = io_cpu_tlb_uncached ? io_cpu_tlb_paddr : _GEN_501; // @[playground/src/cache/ICache.scala 250:41 252:19]
  wire [7:0] _GEN_721 = io_cpu_tlb_uncached ? 8'h0 : _GEN_502; // @[playground/src/cache/ICache.scala 250:41 253:19]
  wire [2:0] _GEN_722 = io_cpu_tlb_uncached ? 3'h2 : _GEN_503; // @[playground/src/cache/ICache.scala 250:41 254:19]
  wire  _GEN_723 = io_cpu_tlb_uncached | _GEN_504; // @[playground/src/cache/ICache.scala 250:41 255:19]
  wire  _GEN_724 = io_cpu_tlb_uncached ? replace_wstrb_0_0_0 : _GEN_505; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_725 = io_cpu_tlb_uncached ? replace_wstrb_1_0_0 : _GEN_506; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_726 = io_cpu_tlb_uncached ? replace_wstrb_0_1_0 : _GEN_507; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_727 = io_cpu_tlb_uncached ? replace_wstrb_1_1_0 : _GEN_508; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_728 = io_cpu_tlb_uncached ? replace_wstrb_0_2_0 : _GEN_509; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_729 = io_cpu_tlb_uncached ? replace_wstrb_1_2_0 : _GEN_510; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_730 = io_cpu_tlb_uncached ? replace_wstrb_0_3_0 : _GEN_511; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_731 = io_cpu_tlb_uncached ? replace_wstrb_1_3_0 : _GEN_512; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_732 = io_cpu_tlb_uncached ? replace_wstrb_0_4_0 : _GEN_513; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_733 = io_cpu_tlb_uncached ? replace_wstrb_1_4_0 : _GEN_514; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_734 = io_cpu_tlb_uncached ? replace_wstrb_0_5_0 : _GEN_515; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_735 = io_cpu_tlb_uncached ? replace_wstrb_1_5_0 : _GEN_516; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_736 = io_cpu_tlb_uncached ? replace_wstrb_0_6_0 : _GEN_517; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_737 = io_cpu_tlb_uncached ? replace_wstrb_1_6_0 : _GEN_518; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_738 = io_cpu_tlb_uncached ? replace_wstrb_0_7_0 : _GEN_519; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_739 = io_cpu_tlb_uncached ? replace_wstrb_1_7_0 : _GEN_520; // @[playground/src/cache/ICache.scala 117:30 250:41]
  wire  _GEN_740 = io_cpu_tlb_uncached ? tag_wstrb_0 : _GEN_521; // @[playground/src/cache/ICache.scala 106:26 250:41]
  wire  _GEN_741 = io_cpu_tlb_uncached ? tag_wstrb_1 : _GEN_522; // @[playground/src/cache/ICache.scala 106:26 250:41]
  wire [19:0] _GEN_742 = io_cpu_tlb_uncached ? tag_wdata : _GEN_523; // @[playground/src/cache/ICache.scala 107:26 250:41]
  wire  _GEN_743 = io_cpu_tlb_uncached ? valid_0_0 : _GEN_524; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_744 = io_cpu_tlb_uncached ? valid_0_1 : _GEN_525; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_745 = io_cpu_tlb_uncached ? valid_0_2 : _GEN_526; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_746 = io_cpu_tlb_uncached ? valid_0_3 : _GEN_527; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_747 = io_cpu_tlb_uncached ? valid_0_4 : _GEN_528; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_748 = io_cpu_tlb_uncached ? valid_0_5 : _GEN_529; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_749 = io_cpu_tlb_uncached ? valid_0_6 : _GEN_530; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_750 = io_cpu_tlb_uncached ? valid_0_7 : _GEN_531; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_751 = io_cpu_tlb_uncached ? valid_0_8 : _GEN_532; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_752 = io_cpu_tlb_uncached ? valid_0_9 : _GEN_533; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_753 = io_cpu_tlb_uncached ? valid_0_10 : _GEN_534; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_754 = io_cpu_tlb_uncached ? valid_0_11 : _GEN_535; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_755 = io_cpu_tlb_uncached ? valid_0_12 : _GEN_536; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_756 = io_cpu_tlb_uncached ? valid_0_13 : _GEN_537; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_757 = io_cpu_tlb_uncached ? valid_0_14 : _GEN_538; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_758 = io_cpu_tlb_uncached ? valid_0_15 : _GEN_539; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_759 = io_cpu_tlb_uncached ? valid_0_16 : _GEN_540; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_760 = io_cpu_tlb_uncached ? valid_0_17 : _GEN_541; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_761 = io_cpu_tlb_uncached ? valid_0_18 : _GEN_542; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_762 = io_cpu_tlb_uncached ? valid_0_19 : _GEN_543; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_763 = io_cpu_tlb_uncached ? valid_0_20 : _GEN_544; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_764 = io_cpu_tlb_uncached ? valid_0_21 : _GEN_545; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_765 = io_cpu_tlb_uncached ? valid_0_22 : _GEN_546; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_766 = io_cpu_tlb_uncached ? valid_0_23 : _GEN_547; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_767 = io_cpu_tlb_uncached ? valid_0_24 : _GEN_548; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_768 = io_cpu_tlb_uncached ? valid_0_25 : _GEN_549; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_769 = io_cpu_tlb_uncached ? valid_0_26 : _GEN_550; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_770 = io_cpu_tlb_uncached ? valid_0_27 : _GEN_551; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_771 = io_cpu_tlb_uncached ? valid_0_28 : _GEN_552; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_772 = io_cpu_tlb_uncached ? valid_0_29 : _GEN_553; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_773 = io_cpu_tlb_uncached ? valid_0_30 : _GEN_554; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_774 = io_cpu_tlb_uncached ? valid_0_31 : _GEN_555; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_775 = io_cpu_tlb_uncached ? valid_0_32 : _GEN_556; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_776 = io_cpu_tlb_uncached ? valid_0_33 : _GEN_557; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_777 = io_cpu_tlb_uncached ? valid_0_34 : _GEN_558; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_778 = io_cpu_tlb_uncached ? valid_0_35 : _GEN_559; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_779 = io_cpu_tlb_uncached ? valid_0_36 : _GEN_560; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_780 = io_cpu_tlb_uncached ? valid_0_37 : _GEN_561; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_781 = io_cpu_tlb_uncached ? valid_0_38 : _GEN_562; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_782 = io_cpu_tlb_uncached ? valid_0_39 : _GEN_563; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_783 = io_cpu_tlb_uncached ? valid_0_40 : _GEN_564; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_784 = io_cpu_tlb_uncached ? valid_0_41 : _GEN_565; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_785 = io_cpu_tlb_uncached ? valid_0_42 : _GEN_566; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_786 = io_cpu_tlb_uncached ? valid_0_43 : _GEN_567; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_787 = io_cpu_tlb_uncached ? valid_0_44 : _GEN_568; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_788 = io_cpu_tlb_uncached ? valid_0_45 : _GEN_569; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_789 = io_cpu_tlb_uncached ? valid_0_46 : _GEN_570; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_790 = io_cpu_tlb_uncached ? valid_0_47 : _GEN_571; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_791 = io_cpu_tlb_uncached ? valid_0_48 : _GEN_572; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_792 = io_cpu_tlb_uncached ? valid_0_49 : _GEN_573; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_793 = io_cpu_tlb_uncached ? valid_0_50 : _GEN_574; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_794 = io_cpu_tlb_uncached ? valid_0_51 : _GEN_575; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_795 = io_cpu_tlb_uncached ? valid_0_52 : _GEN_576; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_796 = io_cpu_tlb_uncached ? valid_0_53 : _GEN_577; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_797 = io_cpu_tlb_uncached ? valid_0_54 : _GEN_578; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_798 = io_cpu_tlb_uncached ? valid_0_55 : _GEN_579; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_799 = io_cpu_tlb_uncached ? valid_0_56 : _GEN_580; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_800 = io_cpu_tlb_uncached ? valid_0_57 : _GEN_581; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_801 = io_cpu_tlb_uncached ? valid_0_58 : _GEN_582; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_802 = io_cpu_tlb_uncached ? valid_0_59 : _GEN_583; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_803 = io_cpu_tlb_uncached ? valid_0_60 : _GEN_584; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_804 = io_cpu_tlb_uncached ? valid_0_61 : _GEN_585; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_805 = io_cpu_tlb_uncached ? valid_0_62 : _GEN_586; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_806 = io_cpu_tlb_uncached ? valid_0_63 : _GEN_587; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_807 = io_cpu_tlb_uncached ? valid_1_0 : _GEN_588; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_808 = io_cpu_tlb_uncached ? valid_1_1 : _GEN_589; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_809 = io_cpu_tlb_uncached ? valid_1_2 : _GEN_590; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_810 = io_cpu_tlb_uncached ? valid_1_3 : _GEN_591; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_811 = io_cpu_tlb_uncached ? valid_1_4 : _GEN_592; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_812 = io_cpu_tlb_uncached ? valid_1_5 : _GEN_593; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_813 = io_cpu_tlb_uncached ? valid_1_6 : _GEN_594; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_814 = io_cpu_tlb_uncached ? valid_1_7 : _GEN_595; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_815 = io_cpu_tlb_uncached ? valid_1_8 : _GEN_596; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_816 = io_cpu_tlb_uncached ? valid_1_9 : _GEN_597; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_817 = io_cpu_tlb_uncached ? valid_1_10 : _GEN_598; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_818 = io_cpu_tlb_uncached ? valid_1_11 : _GEN_599; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_819 = io_cpu_tlb_uncached ? valid_1_12 : _GEN_600; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_820 = io_cpu_tlb_uncached ? valid_1_13 : _GEN_601; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_821 = io_cpu_tlb_uncached ? valid_1_14 : _GEN_602; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_822 = io_cpu_tlb_uncached ? valid_1_15 : _GEN_603; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_823 = io_cpu_tlb_uncached ? valid_1_16 : _GEN_604; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_824 = io_cpu_tlb_uncached ? valid_1_17 : _GEN_605; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_825 = io_cpu_tlb_uncached ? valid_1_18 : _GEN_606; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_826 = io_cpu_tlb_uncached ? valid_1_19 : _GEN_607; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_827 = io_cpu_tlb_uncached ? valid_1_20 : _GEN_608; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_828 = io_cpu_tlb_uncached ? valid_1_21 : _GEN_609; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_829 = io_cpu_tlb_uncached ? valid_1_22 : _GEN_610; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_830 = io_cpu_tlb_uncached ? valid_1_23 : _GEN_611; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_831 = io_cpu_tlb_uncached ? valid_1_24 : _GEN_612; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_832 = io_cpu_tlb_uncached ? valid_1_25 : _GEN_613; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_833 = io_cpu_tlb_uncached ? valid_1_26 : _GEN_614; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_834 = io_cpu_tlb_uncached ? valid_1_27 : _GEN_615; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_835 = io_cpu_tlb_uncached ? valid_1_28 : _GEN_616; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_836 = io_cpu_tlb_uncached ? valid_1_29 : _GEN_617; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_837 = io_cpu_tlb_uncached ? valid_1_30 : _GEN_618; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_838 = io_cpu_tlb_uncached ? valid_1_31 : _GEN_619; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_839 = io_cpu_tlb_uncached ? valid_1_32 : _GEN_620; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_840 = io_cpu_tlb_uncached ? valid_1_33 : _GEN_621; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_841 = io_cpu_tlb_uncached ? valid_1_34 : _GEN_622; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_842 = io_cpu_tlb_uncached ? valid_1_35 : _GEN_623; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_843 = io_cpu_tlb_uncached ? valid_1_36 : _GEN_624; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_844 = io_cpu_tlb_uncached ? valid_1_37 : _GEN_625; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_845 = io_cpu_tlb_uncached ? valid_1_38 : _GEN_626; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_846 = io_cpu_tlb_uncached ? valid_1_39 : _GEN_627; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_847 = io_cpu_tlb_uncached ? valid_1_40 : _GEN_628; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_848 = io_cpu_tlb_uncached ? valid_1_41 : _GEN_629; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_849 = io_cpu_tlb_uncached ? valid_1_42 : _GEN_630; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_850 = io_cpu_tlb_uncached ? valid_1_43 : _GEN_631; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_851 = io_cpu_tlb_uncached ? valid_1_44 : _GEN_632; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_852 = io_cpu_tlb_uncached ? valid_1_45 : _GEN_633; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_853 = io_cpu_tlb_uncached ? valid_1_46 : _GEN_634; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_854 = io_cpu_tlb_uncached ? valid_1_47 : _GEN_635; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_855 = io_cpu_tlb_uncached ? valid_1_48 : _GEN_636; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_856 = io_cpu_tlb_uncached ? valid_1_49 : _GEN_637; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_857 = io_cpu_tlb_uncached ? valid_1_50 : _GEN_638; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_858 = io_cpu_tlb_uncached ? valid_1_51 : _GEN_639; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_859 = io_cpu_tlb_uncached ? valid_1_52 : _GEN_640; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_860 = io_cpu_tlb_uncached ? valid_1_53 : _GEN_641; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_861 = io_cpu_tlb_uncached ? valid_1_54 : _GEN_642; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_862 = io_cpu_tlb_uncached ? valid_1_55 : _GEN_643; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_863 = io_cpu_tlb_uncached ? valid_1_56 : _GEN_644; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_864 = io_cpu_tlb_uncached ? valid_1_57 : _GEN_645; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_865 = io_cpu_tlb_uncached ? valid_1_58 : _GEN_646; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_866 = io_cpu_tlb_uncached ? valid_1_59 : _GEN_647; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_867 = io_cpu_tlb_uncached ? valid_1_60 : _GEN_648; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_868 = io_cpu_tlb_uncached ? valid_1_61 : _GEN_649; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_869 = io_cpu_tlb_uncached ? valid_1_62 : _GEN_650; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_870 = io_cpu_tlb_uncached ? valid_1_63 : _GEN_651; // @[playground/src/cache/ICache.scala 250:41 95:22]
  wire  _GEN_871 = io_cpu_tlb_uncached ? lru_0 : _GEN_652; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_872 = io_cpu_tlb_uncached ? lru_1 : _GEN_653; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_873 = io_cpu_tlb_uncached ? lru_2 : _GEN_654; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_874 = io_cpu_tlb_uncached ? lru_3 : _GEN_655; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_875 = io_cpu_tlb_uncached ? lru_4 : _GEN_656; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_876 = io_cpu_tlb_uncached ? lru_5 : _GEN_657; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_877 = io_cpu_tlb_uncached ? lru_6 : _GEN_658; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_878 = io_cpu_tlb_uncached ? lru_7 : _GEN_659; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_879 = io_cpu_tlb_uncached ? lru_8 : _GEN_660; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_880 = io_cpu_tlb_uncached ? lru_9 : _GEN_661; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_881 = io_cpu_tlb_uncached ? lru_10 : _GEN_662; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_882 = io_cpu_tlb_uncached ? lru_11 : _GEN_663; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_883 = io_cpu_tlb_uncached ? lru_12 : _GEN_664; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_884 = io_cpu_tlb_uncached ? lru_13 : _GEN_665; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_885 = io_cpu_tlb_uncached ? lru_14 : _GEN_666; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_886 = io_cpu_tlb_uncached ? lru_15 : _GEN_667; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_887 = io_cpu_tlb_uncached ? lru_16 : _GEN_668; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_888 = io_cpu_tlb_uncached ? lru_17 : _GEN_669; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_889 = io_cpu_tlb_uncached ? lru_18 : _GEN_670; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_890 = io_cpu_tlb_uncached ? lru_19 : _GEN_671; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_891 = io_cpu_tlb_uncached ? lru_20 : _GEN_672; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_892 = io_cpu_tlb_uncached ? lru_21 : _GEN_673; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_893 = io_cpu_tlb_uncached ? lru_22 : _GEN_674; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_894 = io_cpu_tlb_uncached ? lru_23 : _GEN_675; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_895 = io_cpu_tlb_uncached ? lru_24 : _GEN_676; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_896 = io_cpu_tlb_uncached ? lru_25 : _GEN_677; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_897 = io_cpu_tlb_uncached ? lru_26 : _GEN_678; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_898 = io_cpu_tlb_uncached ? lru_27 : _GEN_679; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_899 = io_cpu_tlb_uncached ? lru_28 : _GEN_680; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_900 = io_cpu_tlb_uncached ? lru_29 : _GEN_681; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_901 = io_cpu_tlb_uncached ? lru_30 : _GEN_682; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_902 = io_cpu_tlb_uncached ? lru_31 : _GEN_683; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_903 = io_cpu_tlb_uncached ? lru_32 : _GEN_684; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_904 = io_cpu_tlb_uncached ? lru_33 : _GEN_685; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_905 = io_cpu_tlb_uncached ? lru_34 : _GEN_686; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_906 = io_cpu_tlb_uncached ? lru_35 : _GEN_687; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_907 = io_cpu_tlb_uncached ? lru_36 : _GEN_688; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_908 = io_cpu_tlb_uncached ? lru_37 : _GEN_689; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_909 = io_cpu_tlb_uncached ? lru_38 : _GEN_690; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_910 = io_cpu_tlb_uncached ? lru_39 : _GEN_691; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_911 = io_cpu_tlb_uncached ? lru_40 : _GEN_692; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_912 = io_cpu_tlb_uncached ? lru_41 : _GEN_693; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_913 = io_cpu_tlb_uncached ? lru_42 : _GEN_694; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_914 = io_cpu_tlb_uncached ? lru_43 : _GEN_695; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_915 = io_cpu_tlb_uncached ? lru_44 : _GEN_696; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_916 = io_cpu_tlb_uncached ? lru_45 : _GEN_697; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_917 = io_cpu_tlb_uncached ? lru_46 : _GEN_698; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_918 = io_cpu_tlb_uncached ? lru_47 : _GEN_699; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_919 = io_cpu_tlb_uncached ? lru_48 : _GEN_700; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_920 = io_cpu_tlb_uncached ? lru_49 : _GEN_701; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_921 = io_cpu_tlb_uncached ? lru_50 : _GEN_702; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_922 = io_cpu_tlb_uncached ? lru_51 : _GEN_703; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_923 = io_cpu_tlb_uncached ? lru_52 : _GEN_704; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_924 = io_cpu_tlb_uncached ? lru_53 : _GEN_705; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_925 = io_cpu_tlb_uncached ? lru_54 : _GEN_706; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_926 = io_cpu_tlb_uncached ? lru_55 : _GEN_707; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_927 = io_cpu_tlb_uncached ? lru_56 : _GEN_708; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_928 = io_cpu_tlb_uncached ? lru_57 : _GEN_709; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_929 = io_cpu_tlb_uncached ? lru_58 : _GEN_710; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_930 = io_cpu_tlb_uncached ? lru_59 : _GEN_711; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_931 = io_cpu_tlb_uncached ? lru_60 : _GEN_712; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_932 = io_cpu_tlb_uncached ? lru_61 : _GEN_713; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_933 = io_cpu_tlb_uncached ? lru_62 : _GEN_714; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire  _GEN_934 = io_cpu_tlb_uncached ? lru_63 : _GEN_715; // @[playground/src/cache/ICache.scala 110:20 250:41]
  wire [31:0] _GEN_935 = io_cpu_tlb_uncached ? rdata_in_wait_1_inst : _GEN_716; // @[playground/src/cache/ICache.scala 149:30 250:41]
  wire  _GEN_936 = io_cpu_tlb_uncached ? rdata_in_wait_0_valid : _GEN_717; // @[playground/src/cache/ICache.scala 149:30 250:41]
  wire  _GEN_937 = io_cpu_tlb_uncached ? rdata_in_wait_1_valid : _GEN_718; // @[playground/src/cache/ICache.scala 149:30 250:41]
  wire [2:0] _GEN_938 = ~io_cpu_tlb_hit ? 3'h5 : _GEN_719; // @[playground/src/cache/ICache.scala 248:37 249:17]
  wire [31:0] _GEN_939 = ~io_cpu_tlb_hit ? ar_addr : _GEN_720; // @[playground/src/cache/ICache.scala 207:24 248:37]
  wire [7:0] _GEN_940 = ~io_cpu_tlb_hit ? ar_len : _GEN_721; // @[playground/src/cache/ICache.scala 207:24 248:37]
  wire [2:0] _GEN_941 = ~io_cpu_tlb_hit ? ar_size : _GEN_722; // @[playground/src/cache/ICache.scala 207:24 248:37]
  wire  _GEN_942 = ~io_cpu_tlb_hit ? arvalid : _GEN_723; // @[playground/src/cache/ICache.scala 208:24 248:37]
  wire  _GEN_943 = ~io_cpu_tlb_hit ? replace_wstrb_0_0_0 : _GEN_724; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_944 = ~io_cpu_tlb_hit ? replace_wstrb_1_0_0 : _GEN_725; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_945 = ~io_cpu_tlb_hit ? replace_wstrb_0_1_0 : _GEN_726; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_946 = ~io_cpu_tlb_hit ? replace_wstrb_1_1_0 : _GEN_727; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_947 = ~io_cpu_tlb_hit ? replace_wstrb_0_2_0 : _GEN_728; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_948 = ~io_cpu_tlb_hit ? replace_wstrb_1_2_0 : _GEN_729; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_949 = ~io_cpu_tlb_hit ? replace_wstrb_0_3_0 : _GEN_730; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_950 = ~io_cpu_tlb_hit ? replace_wstrb_1_3_0 : _GEN_731; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_951 = ~io_cpu_tlb_hit ? replace_wstrb_0_4_0 : _GEN_732; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_952 = ~io_cpu_tlb_hit ? replace_wstrb_1_4_0 : _GEN_733; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_953 = ~io_cpu_tlb_hit ? replace_wstrb_0_5_0 : _GEN_734; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_954 = ~io_cpu_tlb_hit ? replace_wstrb_1_5_0 : _GEN_735; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_955 = ~io_cpu_tlb_hit ? replace_wstrb_0_6_0 : _GEN_736; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_956 = ~io_cpu_tlb_hit ? replace_wstrb_1_6_0 : _GEN_737; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_957 = ~io_cpu_tlb_hit ? replace_wstrb_0_7_0 : _GEN_738; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_958 = ~io_cpu_tlb_hit ? replace_wstrb_1_7_0 : _GEN_739; // @[playground/src/cache/ICache.scala 117:30 248:37]
  wire  _GEN_959 = ~io_cpu_tlb_hit ? tag_wstrb_0 : _GEN_740; // @[playground/src/cache/ICache.scala 106:26 248:37]
  wire  _GEN_960 = ~io_cpu_tlb_hit ? tag_wstrb_1 : _GEN_741; // @[playground/src/cache/ICache.scala 106:26 248:37]
  wire [19:0] _GEN_961 = ~io_cpu_tlb_hit ? tag_wdata : _GEN_742; // @[playground/src/cache/ICache.scala 107:26 248:37]
  wire  _GEN_962 = ~io_cpu_tlb_hit ? valid_0_0 : _GEN_743; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_963 = ~io_cpu_tlb_hit ? valid_0_1 : _GEN_744; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_964 = ~io_cpu_tlb_hit ? valid_0_2 : _GEN_745; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_965 = ~io_cpu_tlb_hit ? valid_0_3 : _GEN_746; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_966 = ~io_cpu_tlb_hit ? valid_0_4 : _GEN_747; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_967 = ~io_cpu_tlb_hit ? valid_0_5 : _GEN_748; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_968 = ~io_cpu_tlb_hit ? valid_0_6 : _GEN_749; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_969 = ~io_cpu_tlb_hit ? valid_0_7 : _GEN_750; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_970 = ~io_cpu_tlb_hit ? valid_0_8 : _GEN_751; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_971 = ~io_cpu_tlb_hit ? valid_0_9 : _GEN_752; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_972 = ~io_cpu_tlb_hit ? valid_0_10 : _GEN_753; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_973 = ~io_cpu_tlb_hit ? valid_0_11 : _GEN_754; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_974 = ~io_cpu_tlb_hit ? valid_0_12 : _GEN_755; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_975 = ~io_cpu_tlb_hit ? valid_0_13 : _GEN_756; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_976 = ~io_cpu_tlb_hit ? valid_0_14 : _GEN_757; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_977 = ~io_cpu_tlb_hit ? valid_0_15 : _GEN_758; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_978 = ~io_cpu_tlb_hit ? valid_0_16 : _GEN_759; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_979 = ~io_cpu_tlb_hit ? valid_0_17 : _GEN_760; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_980 = ~io_cpu_tlb_hit ? valid_0_18 : _GEN_761; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_981 = ~io_cpu_tlb_hit ? valid_0_19 : _GEN_762; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_982 = ~io_cpu_tlb_hit ? valid_0_20 : _GEN_763; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_983 = ~io_cpu_tlb_hit ? valid_0_21 : _GEN_764; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_984 = ~io_cpu_tlb_hit ? valid_0_22 : _GEN_765; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_985 = ~io_cpu_tlb_hit ? valid_0_23 : _GEN_766; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_986 = ~io_cpu_tlb_hit ? valid_0_24 : _GEN_767; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_987 = ~io_cpu_tlb_hit ? valid_0_25 : _GEN_768; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_988 = ~io_cpu_tlb_hit ? valid_0_26 : _GEN_769; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_989 = ~io_cpu_tlb_hit ? valid_0_27 : _GEN_770; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_990 = ~io_cpu_tlb_hit ? valid_0_28 : _GEN_771; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_991 = ~io_cpu_tlb_hit ? valid_0_29 : _GEN_772; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_992 = ~io_cpu_tlb_hit ? valid_0_30 : _GEN_773; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_993 = ~io_cpu_tlb_hit ? valid_0_31 : _GEN_774; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_994 = ~io_cpu_tlb_hit ? valid_0_32 : _GEN_775; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_995 = ~io_cpu_tlb_hit ? valid_0_33 : _GEN_776; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_996 = ~io_cpu_tlb_hit ? valid_0_34 : _GEN_777; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_997 = ~io_cpu_tlb_hit ? valid_0_35 : _GEN_778; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_998 = ~io_cpu_tlb_hit ? valid_0_36 : _GEN_779; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_999 = ~io_cpu_tlb_hit ? valid_0_37 : _GEN_780; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1000 = ~io_cpu_tlb_hit ? valid_0_38 : _GEN_781; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1001 = ~io_cpu_tlb_hit ? valid_0_39 : _GEN_782; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1002 = ~io_cpu_tlb_hit ? valid_0_40 : _GEN_783; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1003 = ~io_cpu_tlb_hit ? valid_0_41 : _GEN_784; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1004 = ~io_cpu_tlb_hit ? valid_0_42 : _GEN_785; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1005 = ~io_cpu_tlb_hit ? valid_0_43 : _GEN_786; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1006 = ~io_cpu_tlb_hit ? valid_0_44 : _GEN_787; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1007 = ~io_cpu_tlb_hit ? valid_0_45 : _GEN_788; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1008 = ~io_cpu_tlb_hit ? valid_0_46 : _GEN_789; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1009 = ~io_cpu_tlb_hit ? valid_0_47 : _GEN_790; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1010 = ~io_cpu_tlb_hit ? valid_0_48 : _GEN_791; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1011 = ~io_cpu_tlb_hit ? valid_0_49 : _GEN_792; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1012 = ~io_cpu_tlb_hit ? valid_0_50 : _GEN_793; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1013 = ~io_cpu_tlb_hit ? valid_0_51 : _GEN_794; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1014 = ~io_cpu_tlb_hit ? valid_0_52 : _GEN_795; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1015 = ~io_cpu_tlb_hit ? valid_0_53 : _GEN_796; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1016 = ~io_cpu_tlb_hit ? valid_0_54 : _GEN_797; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1017 = ~io_cpu_tlb_hit ? valid_0_55 : _GEN_798; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1018 = ~io_cpu_tlb_hit ? valid_0_56 : _GEN_799; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1019 = ~io_cpu_tlb_hit ? valid_0_57 : _GEN_800; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1020 = ~io_cpu_tlb_hit ? valid_0_58 : _GEN_801; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1021 = ~io_cpu_tlb_hit ? valid_0_59 : _GEN_802; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1022 = ~io_cpu_tlb_hit ? valid_0_60 : _GEN_803; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1023 = ~io_cpu_tlb_hit ? valid_0_61 : _GEN_804; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1024 = ~io_cpu_tlb_hit ? valid_0_62 : _GEN_805; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1025 = ~io_cpu_tlb_hit ? valid_0_63 : _GEN_806; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1026 = ~io_cpu_tlb_hit ? valid_1_0 : _GEN_807; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1027 = ~io_cpu_tlb_hit ? valid_1_1 : _GEN_808; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1028 = ~io_cpu_tlb_hit ? valid_1_2 : _GEN_809; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1029 = ~io_cpu_tlb_hit ? valid_1_3 : _GEN_810; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1030 = ~io_cpu_tlb_hit ? valid_1_4 : _GEN_811; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1031 = ~io_cpu_tlb_hit ? valid_1_5 : _GEN_812; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1032 = ~io_cpu_tlb_hit ? valid_1_6 : _GEN_813; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1033 = ~io_cpu_tlb_hit ? valid_1_7 : _GEN_814; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1034 = ~io_cpu_tlb_hit ? valid_1_8 : _GEN_815; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1035 = ~io_cpu_tlb_hit ? valid_1_9 : _GEN_816; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1036 = ~io_cpu_tlb_hit ? valid_1_10 : _GEN_817; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1037 = ~io_cpu_tlb_hit ? valid_1_11 : _GEN_818; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1038 = ~io_cpu_tlb_hit ? valid_1_12 : _GEN_819; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1039 = ~io_cpu_tlb_hit ? valid_1_13 : _GEN_820; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1040 = ~io_cpu_tlb_hit ? valid_1_14 : _GEN_821; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1041 = ~io_cpu_tlb_hit ? valid_1_15 : _GEN_822; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1042 = ~io_cpu_tlb_hit ? valid_1_16 : _GEN_823; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1043 = ~io_cpu_tlb_hit ? valid_1_17 : _GEN_824; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1044 = ~io_cpu_tlb_hit ? valid_1_18 : _GEN_825; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1045 = ~io_cpu_tlb_hit ? valid_1_19 : _GEN_826; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1046 = ~io_cpu_tlb_hit ? valid_1_20 : _GEN_827; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1047 = ~io_cpu_tlb_hit ? valid_1_21 : _GEN_828; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1048 = ~io_cpu_tlb_hit ? valid_1_22 : _GEN_829; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1049 = ~io_cpu_tlb_hit ? valid_1_23 : _GEN_830; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1050 = ~io_cpu_tlb_hit ? valid_1_24 : _GEN_831; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1051 = ~io_cpu_tlb_hit ? valid_1_25 : _GEN_832; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1052 = ~io_cpu_tlb_hit ? valid_1_26 : _GEN_833; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1053 = ~io_cpu_tlb_hit ? valid_1_27 : _GEN_834; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1054 = ~io_cpu_tlb_hit ? valid_1_28 : _GEN_835; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1055 = ~io_cpu_tlb_hit ? valid_1_29 : _GEN_836; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1056 = ~io_cpu_tlb_hit ? valid_1_30 : _GEN_837; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1057 = ~io_cpu_tlb_hit ? valid_1_31 : _GEN_838; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1058 = ~io_cpu_tlb_hit ? valid_1_32 : _GEN_839; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1059 = ~io_cpu_tlb_hit ? valid_1_33 : _GEN_840; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1060 = ~io_cpu_tlb_hit ? valid_1_34 : _GEN_841; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1061 = ~io_cpu_tlb_hit ? valid_1_35 : _GEN_842; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1062 = ~io_cpu_tlb_hit ? valid_1_36 : _GEN_843; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1063 = ~io_cpu_tlb_hit ? valid_1_37 : _GEN_844; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1064 = ~io_cpu_tlb_hit ? valid_1_38 : _GEN_845; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1065 = ~io_cpu_tlb_hit ? valid_1_39 : _GEN_846; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1066 = ~io_cpu_tlb_hit ? valid_1_40 : _GEN_847; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1067 = ~io_cpu_tlb_hit ? valid_1_41 : _GEN_848; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1068 = ~io_cpu_tlb_hit ? valid_1_42 : _GEN_849; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1069 = ~io_cpu_tlb_hit ? valid_1_43 : _GEN_850; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1070 = ~io_cpu_tlb_hit ? valid_1_44 : _GEN_851; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1071 = ~io_cpu_tlb_hit ? valid_1_45 : _GEN_852; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1072 = ~io_cpu_tlb_hit ? valid_1_46 : _GEN_853; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1073 = ~io_cpu_tlb_hit ? valid_1_47 : _GEN_854; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1074 = ~io_cpu_tlb_hit ? valid_1_48 : _GEN_855; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1075 = ~io_cpu_tlb_hit ? valid_1_49 : _GEN_856; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1076 = ~io_cpu_tlb_hit ? valid_1_50 : _GEN_857; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1077 = ~io_cpu_tlb_hit ? valid_1_51 : _GEN_858; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1078 = ~io_cpu_tlb_hit ? valid_1_52 : _GEN_859; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1079 = ~io_cpu_tlb_hit ? valid_1_53 : _GEN_860; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1080 = ~io_cpu_tlb_hit ? valid_1_54 : _GEN_861; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1081 = ~io_cpu_tlb_hit ? valid_1_55 : _GEN_862; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1082 = ~io_cpu_tlb_hit ? valid_1_56 : _GEN_863; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1083 = ~io_cpu_tlb_hit ? valid_1_57 : _GEN_864; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1084 = ~io_cpu_tlb_hit ? valid_1_58 : _GEN_865; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1085 = ~io_cpu_tlb_hit ? valid_1_59 : _GEN_866; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1086 = ~io_cpu_tlb_hit ? valid_1_60 : _GEN_867; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1087 = ~io_cpu_tlb_hit ? valid_1_61 : _GEN_868; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1088 = ~io_cpu_tlb_hit ? valid_1_62 : _GEN_869; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1089 = ~io_cpu_tlb_hit ? valid_1_63 : _GEN_870; // @[playground/src/cache/ICache.scala 248:37 95:22]
  wire  _GEN_1090 = ~io_cpu_tlb_hit ? lru_0 : _GEN_871; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1091 = ~io_cpu_tlb_hit ? lru_1 : _GEN_872; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1092 = ~io_cpu_tlb_hit ? lru_2 : _GEN_873; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1093 = ~io_cpu_tlb_hit ? lru_3 : _GEN_874; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1094 = ~io_cpu_tlb_hit ? lru_4 : _GEN_875; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1095 = ~io_cpu_tlb_hit ? lru_5 : _GEN_876; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1096 = ~io_cpu_tlb_hit ? lru_6 : _GEN_877; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1097 = ~io_cpu_tlb_hit ? lru_7 : _GEN_878; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1098 = ~io_cpu_tlb_hit ? lru_8 : _GEN_879; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1099 = ~io_cpu_tlb_hit ? lru_9 : _GEN_880; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1100 = ~io_cpu_tlb_hit ? lru_10 : _GEN_881; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1101 = ~io_cpu_tlb_hit ? lru_11 : _GEN_882; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1102 = ~io_cpu_tlb_hit ? lru_12 : _GEN_883; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1103 = ~io_cpu_tlb_hit ? lru_13 : _GEN_884; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1104 = ~io_cpu_tlb_hit ? lru_14 : _GEN_885; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1105 = ~io_cpu_tlb_hit ? lru_15 : _GEN_886; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1106 = ~io_cpu_tlb_hit ? lru_16 : _GEN_887; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1107 = ~io_cpu_tlb_hit ? lru_17 : _GEN_888; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1108 = ~io_cpu_tlb_hit ? lru_18 : _GEN_889; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1109 = ~io_cpu_tlb_hit ? lru_19 : _GEN_890; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1110 = ~io_cpu_tlb_hit ? lru_20 : _GEN_891; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1111 = ~io_cpu_tlb_hit ? lru_21 : _GEN_892; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1112 = ~io_cpu_tlb_hit ? lru_22 : _GEN_893; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1113 = ~io_cpu_tlb_hit ? lru_23 : _GEN_894; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1114 = ~io_cpu_tlb_hit ? lru_24 : _GEN_895; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1115 = ~io_cpu_tlb_hit ? lru_25 : _GEN_896; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1116 = ~io_cpu_tlb_hit ? lru_26 : _GEN_897; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1117 = ~io_cpu_tlb_hit ? lru_27 : _GEN_898; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1118 = ~io_cpu_tlb_hit ? lru_28 : _GEN_899; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1119 = ~io_cpu_tlb_hit ? lru_29 : _GEN_900; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1120 = ~io_cpu_tlb_hit ? lru_30 : _GEN_901; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1121 = ~io_cpu_tlb_hit ? lru_31 : _GEN_902; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1122 = ~io_cpu_tlb_hit ? lru_32 : _GEN_903; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1123 = ~io_cpu_tlb_hit ? lru_33 : _GEN_904; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1124 = ~io_cpu_tlb_hit ? lru_34 : _GEN_905; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1125 = ~io_cpu_tlb_hit ? lru_35 : _GEN_906; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1126 = ~io_cpu_tlb_hit ? lru_36 : _GEN_907; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1127 = ~io_cpu_tlb_hit ? lru_37 : _GEN_908; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1128 = ~io_cpu_tlb_hit ? lru_38 : _GEN_909; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1129 = ~io_cpu_tlb_hit ? lru_39 : _GEN_910; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1130 = ~io_cpu_tlb_hit ? lru_40 : _GEN_911; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1131 = ~io_cpu_tlb_hit ? lru_41 : _GEN_912; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1132 = ~io_cpu_tlb_hit ? lru_42 : _GEN_913; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1133 = ~io_cpu_tlb_hit ? lru_43 : _GEN_914; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1134 = ~io_cpu_tlb_hit ? lru_44 : _GEN_915; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1135 = ~io_cpu_tlb_hit ? lru_45 : _GEN_916; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1136 = ~io_cpu_tlb_hit ? lru_46 : _GEN_917; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1137 = ~io_cpu_tlb_hit ? lru_47 : _GEN_918; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1138 = ~io_cpu_tlb_hit ? lru_48 : _GEN_919; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1139 = ~io_cpu_tlb_hit ? lru_49 : _GEN_920; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1140 = ~io_cpu_tlb_hit ? lru_50 : _GEN_921; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1141 = ~io_cpu_tlb_hit ? lru_51 : _GEN_922; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1142 = ~io_cpu_tlb_hit ? lru_52 : _GEN_923; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1143 = ~io_cpu_tlb_hit ? lru_53 : _GEN_924; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1144 = ~io_cpu_tlb_hit ? lru_54 : _GEN_925; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1145 = ~io_cpu_tlb_hit ? lru_55 : _GEN_926; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1146 = ~io_cpu_tlb_hit ? lru_56 : _GEN_927; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1147 = ~io_cpu_tlb_hit ? lru_57 : _GEN_928; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1148 = ~io_cpu_tlb_hit ? lru_58 : _GEN_929; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1149 = ~io_cpu_tlb_hit ? lru_59 : _GEN_930; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1150 = ~io_cpu_tlb_hit ? lru_60 : _GEN_931; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1151 = ~io_cpu_tlb_hit ? lru_61 : _GEN_932; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1152 = ~io_cpu_tlb_hit ? lru_62 : _GEN_933; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire  _GEN_1153 = ~io_cpu_tlb_hit ? lru_63 : _GEN_934; // @[playground/src/cache/ICache.scala 110:20 248:37]
  wire [31:0] _GEN_1154 = ~io_cpu_tlb_hit ? rdata_in_wait_1_inst : _GEN_935; // @[playground/src/cache/ICache.scala 149:30 248:37]
  wire  _GEN_1155 = ~io_cpu_tlb_hit ? rdata_in_wait_0_valid : _GEN_936; // @[playground/src/cache/ICache.scala 149:30 248:37]
  wire  _GEN_1156 = ~io_cpu_tlb_hit ? rdata_in_wait_1_valid : _GEN_937; // @[playground/src/cache/ICache.scala 149:30 248:37]
  wire  _GEN_1157 = addr_err & _addr_err_T_101; // @[playground/src/cache/ICache.scala 237:23 239:24]
  wire  _GEN_1158 = addr_err & _GEN_151; // @[playground/src/cache/ICache.scala 235:23 239:24]
  wire [2:0] _GEN_1159 = addr_err ? 3'h3 : _GEN_938; // @[playground/src/cache/ICache.scala 239:24 245:34]
  wire  _GEN_1161 = addr_err | _GEN_1155; // @[playground/src/cache/ICache.scala 239:24 247:34]
  wire  _GEN_1185 = addr_err ? valid_0_0 : _GEN_962; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1186 = addr_err ? valid_0_1 : _GEN_963; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1187 = addr_err ? valid_0_2 : _GEN_964; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1188 = addr_err ? valid_0_3 : _GEN_965; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1189 = addr_err ? valid_0_4 : _GEN_966; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1190 = addr_err ? valid_0_5 : _GEN_967; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1191 = addr_err ? valid_0_6 : _GEN_968; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1192 = addr_err ? valid_0_7 : _GEN_969; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1193 = addr_err ? valid_0_8 : _GEN_970; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1194 = addr_err ? valid_0_9 : _GEN_971; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1195 = addr_err ? valid_0_10 : _GEN_972; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1196 = addr_err ? valid_0_11 : _GEN_973; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1197 = addr_err ? valid_0_12 : _GEN_974; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1198 = addr_err ? valid_0_13 : _GEN_975; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1199 = addr_err ? valid_0_14 : _GEN_976; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1200 = addr_err ? valid_0_15 : _GEN_977; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1201 = addr_err ? valid_0_16 : _GEN_978; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1202 = addr_err ? valid_0_17 : _GEN_979; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1203 = addr_err ? valid_0_18 : _GEN_980; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1204 = addr_err ? valid_0_19 : _GEN_981; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1205 = addr_err ? valid_0_20 : _GEN_982; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1206 = addr_err ? valid_0_21 : _GEN_983; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1207 = addr_err ? valid_0_22 : _GEN_984; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1208 = addr_err ? valid_0_23 : _GEN_985; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1209 = addr_err ? valid_0_24 : _GEN_986; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1210 = addr_err ? valid_0_25 : _GEN_987; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1211 = addr_err ? valid_0_26 : _GEN_988; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1212 = addr_err ? valid_0_27 : _GEN_989; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1213 = addr_err ? valid_0_28 : _GEN_990; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1214 = addr_err ? valid_0_29 : _GEN_991; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1215 = addr_err ? valid_0_30 : _GEN_992; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1216 = addr_err ? valid_0_31 : _GEN_993; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1217 = addr_err ? valid_0_32 : _GEN_994; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1218 = addr_err ? valid_0_33 : _GEN_995; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1219 = addr_err ? valid_0_34 : _GEN_996; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1220 = addr_err ? valid_0_35 : _GEN_997; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1221 = addr_err ? valid_0_36 : _GEN_998; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1222 = addr_err ? valid_0_37 : _GEN_999; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1223 = addr_err ? valid_0_38 : _GEN_1000; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1224 = addr_err ? valid_0_39 : _GEN_1001; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1225 = addr_err ? valid_0_40 : _GEN_1002; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1226 = addr_err ? valid_0_41 : _GEN_1003; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1227 = addr_err ? valid_0_42 : _GEN_1004; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1228 = addr_err ? valid_0_43 : _GEN_1005; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1229 = addr_err ? valid_0_44 : _GEN_1006; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1230 = addr_err ? valid_0_45 : _GEN_1007; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1231 = addr_err ? valid_0_46 : _GEN_1008; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1232 = addr_err ? valid_0_47 : _GEN_1009; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1233 = addr_err ? valid_0_48 : _GEN_1010; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1234 = addr_err ? valid_0_49 : _GEN_1011; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1235 = addr_err ? valid_0_50 : _GEN_1012; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1236 = addr_err ? valid_0_51 : _GEN_1013; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1237 = addr_err ? valid_0_52 : _GEN_1014; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1238 = addr_err ? valid_0_53 : _GEN_1015; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1239 = addr_err ? valid_0_54 : _GEN_1016; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1240 = addr_err ? valid_0_55 : _GEN_1017; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1241 = addr_err ? valid_0_56 : _GEN_1018; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1242 = addr_err ? valid_0_57 : _GEN_1019; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1243 = addr_err ? valid_0_58 : _GEN_1020; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1244 = addr_err ? valid_0_59 : _GEN_1021; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1245 = addr_err ? valid_0_60 : _GEN_1022; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1246 = addr_err ? valid_0_61 : _GEN_1023; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1247 = addr_err ? valid_0_62 : _GEN_1024; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1248 = addr_err ? valid_0_63 : _GEN_1025; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1249 = addr_err ? valid_1_0 : _GEN_1026; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1250 = addr_err ? valid_1_1 : _GEN_1027; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1251 = addr_err ? valid_1_2 : _GEN_1028; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1252 = addr_err ? valid_1_3 : _GEN_1029; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1253 = addr_err ? valid_1_4 : _GEN_1030; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1254 = addr_err ? valid_1_5 : _GEN_1031; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1255 = addr_err ? valid_1_6 : _GEN_1032; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1256 = addr_err ? valid_1_7 : _GEN_1033; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1257 = addr_err ? valid_1_8 : _GEN_1034; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1258 = addr_err ? valid_1_9 : _GEN_1035; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1259 = addr_err ? valid_1_10 : _GEN_1036; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1260 = addr_err ? valid_1_11 : _GEN_1037; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1261 = addr_err ? valid_1_12 : _GEN_1038; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1262 = addr_err ? valid_1_13 : _GEN_1039; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1263 = addr_err ? valid_1_14 : _GEN_1040; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1264 = addr_err ? valid_1_15 : _GEN_1041; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1265 = addr_err ? valid_1_16 : _GEN_1042; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1266 = addr_err ? valid_1_17 : _GEN_1043; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1267 = addr_err ? valid_1_18 : _GEN_1044; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1268 = addr_err ? valid_1_19 : _GEN_1045; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1269 = addr_err ? valid_1_20 : _GEN_1046; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1270 = addr_err ? valid_1_21 : _GEN_1047; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1271 = addr_err ? valid_1_22 : _GEN_1048; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1272 = addr_err ? valid_1_23 : _GEN_1049; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1273 = addr_err ? valid_1_24 : _GEN_1050; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1274 = addr_err ? valid_1_25 : _GEN_1051; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1275 = addr_err ? valid_1_26 : _GEN_1052; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1276 = addr_err ? valid_1_27 : _GEN_1053; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1277 = addr_err ? valid_1_28 : _GEN_1054; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1278 = addr_err ? valid_1_29 : _GEN_1055; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1279 = addr_err ? valid_1_30 : _GEN_1056; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1280 = addr_err ? valid_1_31 : _GEN_1057; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1281 = addr_err ? valid_1_32 : _GEN_1058; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1282 = addr_err ? valid_1_33 : _GEN_1059; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1283 = addr_err ? valid_1_34 : _GEN_1060; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1284 = addr_err ? valid_1_35 : _GEN_1061; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1285 = addr_err ? valid_1_36 : _GEN_1062; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1286 = addr_err ? valid_1_37 : _GEN_1063; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1287 = addr_err ? valid_1_38 : _GEN_1064; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1288 = addr_err ? valid_1_39 : _GEN_1065; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1289 = addr_err ? valid_1_40 : _GEN_1066; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1290 = addr_err ? valid_1_41 : _GEN_1067; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1291 = addr_err ? valid_1_42 : _GEN_1068; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1292 = addr_err ? valid_1_43 : _GEN_1069; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1293 = addr_err ? valid_1_44 : _GEN_1070; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1294 = addr_err ? valid_1_45 : _GEN_1071; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1295 = addr_err ? valid_1_46 : _GEN_1072; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1296 = addr_err ? valid_1_47 : _GEN_1073; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1297 = addr_err ? valid_1_48 : _GEN_1074; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1298 = addr_err ? valid_1_49 : _GEN_1075; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1299 = addr_err ? valid_1_50 : _GEN_1076; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1300 = addr_err ? valid_1_51 : _GEN_1077; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1301 = addr_err ? valid_1_52 : _GEN_1078; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1302 = addr_err ? valid_1_53 : _GEN_1079; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1303 = addr_err ? valid_1_54 : _GEN_1080; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1304 = addr_err ? valid_1_55 : _GEN_1081; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1305 = addr_err ? valid_1_56 : _GEN_1082; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1306 = addr_err ? valid_1_57 : _GEN_1083; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1307 = addr_err ? valid_1_58 : _GEN_1084; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1308 = addr_err ? valid_1_59 : _GEN_1085; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1309 = addr_err ? valid_1_60 : _GEN_1086; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1310 = addr_err ? valid_1_61 : _GEN_1087; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1311 = addr_err ? valid_1_62 : _GEN_1088; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1312 = addr_err ? valid_1_63 : _GEN_1089; // @[playground/src/cache/ICache.scala 239:24 95:22]
  wire  _GEN_1379 = io_cpu_req & _GEN_1157; // @[playground/src/cache/ICache.scala 237:23 238:24]
  wire  _GEN_1380 = io_cpu_req & _GEN_1158; // @[playground/src/cache/ICache.scala 235:23 238:24]
  wire  _GEN_1601 = io_axi_ar_ready ? 1'h0 : arvalid; // @[playground/src/cache/ICache.scala 281:31 282:19 208:24]
  wire  _GEN_1602 = io_axi_ar_ready | rready; // @[playground/src/cache/ICache.scala 281:31 283:19 213:23]
  wire  _T_8 = io_axi_r_ready & io_axi_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [31:0] _rdata_in_wait_0_inst_T_3 = ar_addr[2] ? io_axi_r_bits_data[63:32] : io_axi_r_bits_data[31:0]; // @[playground/src/cache/ICache.scala 287:38]
  wire [31:0] _GEN_1603 = _T_8 ? _rdata_in_wait_0_inst_T_3 : rdata_in_wait_0_inst; // @[playground/src/cache/ICache.scala 149:30 285:33 287:32]
  wire  _GEN_1604 = _T_8 | rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 149:30 285:33 288:32]
  wire  _GEN_1605 = _T_8 ? 1'h0 : rready; // @[playground/src/cache/ICache.scala 213:23 285:33 289:32]
  wire  _GEN_1606 = _T_8 ? io_axi_r_bits_resp != 2'h0 : access_fault; // @[playground/src/cache/ICache.scala 217:32 285:33 290:32]
  wire [2:0] _GEN_1607 = _T_8 ? 3'h3 : state; // @[playground/src/cache/ICache.scala 285:33 291:32 92:94]
  wire  _GEN_1608 = io_axi_ar_valid ? _GEN_1601 : arvalid; // @[playground/src/cache/ICache.scala 208:24 280:29]
  wire [2:0] _GEN_1613 = io_axi_ar_valid ? state : _GEN_1607; // @[playground/src/cache/ICache.scala 280:29 92:94]
  wire  _GEN_1615 = _GEN_215 ? replace_wstrb_1_1_0 : replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1617 = _GEN_215 ? replace_wstrb_1_0_0 : replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1619 = _GEN_215 ? replace_wstrb_1_3_0 : replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1621 = _GEN_215 ? replace_wstrb_1_2_0 : replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1623 = _GEN_215 ? replace_wstrb_1_5_0 : replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1625 = _GEN_215 ? replace_wstrb_1_4_0 : replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1627 = _GEN_215 ? replace_wstrb_1_7_0 : replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire  _GEN_1629 = _GEN_215 ? replace_wstrb_1_6_0 : replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 305:{42,42}]
  wire [7:0] _T_12 = {_GEN_1627,_GEN_1629,_GEN_1623,_GEN_1625,_GEN_1619,_GEN_1621,_GEN_1615,_GEN_1617}; // @[playground/src/cache/ICache.scala 305:42]
  wire [8:0] _T_13 = {_T_12, 1'h0}; // @[playground/src/cache/ICache.scala 305:49]
  wire  _GEN_1630 = ~_GEN_215 ? _T_13[0] : replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1631 = _GEN_215 ? _T_13[0] : replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1632 = ~_GEN_215 ? _T_13[1] : replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1633 = _GEN_215 ? _T_13[1] : replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1634 = ~_GEN_215 ? _T_13[2] : replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1635 = _GEN_215 ? _T_13[2] : replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1636 = ~_GEN_215 ? _T_13[3] : replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1637 = _GEN_215 ? _T_13[3] : replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1638 = ~_GEN_215 ? _T_13[4] : replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1639 = _GEN_215 ? _T_13[4] : replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1640 = ~_GEN_215 ? _T_13[5] : replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1641 = _GEN_215 ? _T_13[5] : replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1642 = ~_GEN_215 ? _T_13[6] : replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1643 = _GEN_215 ? _T_13[6] : replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1644 = ~_GEN_215 ? _T_13[7] : replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1645 = _GEN_215 ? _T_13[7] : replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 117:30 304:{38,38}]
  wire  _GEN_1662 = ~_GEN_215 ? 1'h0 : tag_wstrb_0; // @[playground/src/cache/ICache.scala 106:26 309:{34,34}]
  wire  _GEN_1663 = _GEN_215 ? 1'h0 : tag_wstrb_1; // @[playground/src/cache/ICache.scala 106:26 309:{34,34}]
  wire  _GEN_1664 = ~io_axi_r_bits_last ? _GEN_1630 : _GEN_216; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1665 = ~io_axi_r_bits_last ? _GEN_1631 : _GEN_217; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1666 = ~io_axi_r_bits_last ? _GEN_1632 : _GEN_218; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1667 = ~io_axi_r_bits_last ? _GEN_1633 : _GEN_219; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1668 = ~io_axi_r_bits_last ? _GEN_1634 : _GEN_220; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1669 = ~io_axi_r_bits_last ? _GEN_1635 : _GEN_221; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1670 = ~io_axi_r_bits_last ? _GEN_1636 : _GEN_222; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1671 = ~io_axi_r_bits_last ? _GEN_1637 : _GEN_223; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1672 = ~io_axi_r_bits_last ? _GEN_1638 : _GEN_224; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1673 = ~io_axi_r_bits_last ? _GEN_1639 : _GEN_225; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1674 = ~io_axi_r_bits_last ? _GEN_1640 : _GEN_226; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1675 = ~io_axi_r_bits_last ? _GEN_1641 : _GEN_227; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1676 = ~io_axi_r_bits_last ? _GEN_1642 : _GEN_228; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1677 = ~io_axi_r_bits_last ? _GEN_1643 : _GEN_229; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1678 = ~io_axi_r_bits_last ? _GEN_1644 : _GEN_230; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1679 = ~io_axi_r_bits_last ? _GEN_1645 : _GEN_231; // @[playground/src/cache/ICache.scala 302:35]
  wire  _GEN_1680 = ~io_axi_r_bits_last & rready; // @[playground/src/cache/ICache.scala 213:23 302:35 307:18]
  wire  _GEN_1681 = ~io_axi_r_bits_last ? tag_wstrb_0 : _GEN_1662; // @[playground/src/cache/ICache.scala 106:26 302:35]
  wire  _GEN_1682 = ~io_axi_r_bits_last ? tag_wstrb_1 : _GEN_1663; // @[playground/src/cache/ICache.scala 106:26 302:35]
  wire [2:0] _GEN_1683 = ~io_axi_r_ready ? 3'h0 : state; // @[playground/src/cache/ICache.scala 311:35 312:15 92:94]
  wire  _GEN_1684 = _T_8 ? _GEN_1664 : replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1685 = _T_8 ? _GEN_1665 : replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1686 = _T_8 ? _GEN_1666 : replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1687 = _T_8 ? _GEN_1667 : replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1688 = _T_8 ? _GEN_1668 : replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1689 = _T_8 ? _GEN_1669 : replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1690 = _T_8 ? _GEN_1670 : replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1691 = _T_8 ? _GEN_1671 : replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1692 = _T_8 ? _GEN_1672 : replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1693 = _T_8 ? _GEN_1673 : replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1694 = _T_8 ? _GEN_1674 : replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1695 = _T_8 ? _GEN_1675 : replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1696 = _T_8 ? _GEN_1676 : replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1697 = _T_8 ? _GEN_1677 : replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1698 = _T_8 ? _GEN_1678 : replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1699 = _T_8 ? _GEN_1679 : replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 117:30 300:33]
  wire  _GEN_1700 = _T_8 ? _GEN_1680 : rready; // @[playground/src/cache/ICache.scala 213:23 300:33]
  wire  _GEN_1701 = _T_8 ? _GEN_1681 : tag_wstrb_0; // @[playground/src/cache/ICache.scala 106:26 300:33]
  wire  _GEN_1702 = _T_8 ? _GEN_1682 : tag_wstrb_1; // @[playground/src/cache/ICache.scala 106:26 300:33]
  wire [2:0] _GEN_1703 = _T_8 ? state : _GEN_1683; // @[playground/src/cache/ICache.scala 300:33 92:94]
  wire  _GEN_1704 = io_axi_ar_valid ? _GEN_1602 : _GEN_1700; // @[playground/src/cache/ICache.scala 295:29]
  wire  _GEN_1705 = io_axi_ar_valid ? replace_wstrb_0_0_0 : _GEN_1684; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1706 = io_axi_ar_valid ? replace_wstrb_1_0_0 : _GEN_1685; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1707 = io_axi_ar_valid ? replace_wstrb_0_1_0 : _GEN_1686; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1708 = io_axi_ar_valid ? replace_wstrb_1_1_0 : _GEN_1687; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1709 = io_axi_ar_valid ? replace_wstrb_0_2_0 : _GEN_1688; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1710 = io_axi_ar_valid ? replace_wstrb_1_2_0 : _GEN_1689; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1711 = io_axi_ar_valid ? replace_wstrb_0_3_0 : _GEN_1690; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1712 = io_axi_ar_valid ? replace_wstrb_1_3_0 : _GEN_1691; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1713 = io_axi_ar_valid ? replace_wstrb_0_4_0 : _GEN_1692; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1714 = io_axi_ar_valid ? replace_wstrb_1_4_0 : _GEN_1693; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1715 = io_axi_ar_valid ? replace_wstrb_0_5_0 : _GEN_1694; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1716 = io_axi_ar_valid ? replace_wstrb_1_5_0 : _GEN_1695; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1717 = io_axi_ar_valid ? replace_wstrb_0_6_0 : _GEN_1696; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1718 = io_axi_ar_valid ? replace_wstrb_1_6_0 : _GEN_1697; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1719 = io_axi_ar_valid ? replace_wstrb_0_7_0 : _GEN_1698; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1720 = io_axi_ar_valid ? replace_wstrb_1_7_0 : _GEN_1699; // @[playground/src/cache/ICache.scala 295:29 117:30]
  wire  _GEN_1721 = io_axi_ar_valid ? tag_wstrb_0 : _GEN_1701; // @[playground/src/cache/ICache.scala 106:26 295:29]
  wire  _GEN_1722 = io_axi_ar_valid ? tag_wstrb_1 : _GEN_1702; // @[playground/src/cache/ICache.scala 106:26 295:29]
  wire [2:0] _GEN_1723 = io_axi_ar_valid ? state : _GEN_1703; // @[playground/src/cache/ICache.scala 295:29 92:94]
  wire  _GEN_1724 = io_cpu_complete_single_request ? 1'h0 : access_fault; // @[playground/src/cache/ICache.scala 317:44 318:25 217:32]
  wire  _GEN_1725 = io_cpu_complete_single_request ? 1'h0 : page_fault; // @[playground/src/cache/ICache.scala 317:44 319:25 218:32]
  wire  _GEN_1726 = io_cpu_complete_single_request ? 1'h0 : addr_misaligned; // @[playground/src/cache/ICache.scala 317:44 320:25 219:32]
  wire [2:0] _GEN_1727 = io_cpu_complete_single_request ? 3'h0 : state; // @[playground/src/cache/ICache.scala 317:44 321:25 92:94]
  wire  _GEN_1728 = io_cpu_complete_single_request ? 1'h0 : rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 149:30 317:44 322:68]
  wire  _GEN_1729 = io_cpu_complete_single_request ? 1'h0 : rdata_in_wait_1_valid; // @[playground/src/cache/ICache.scala 149:30 317:44 322:68]
  wire [2:0] _GEN_1730 = ~io_cpu_dcache_stall & ~io_axi_r_valid ? 3'h0 : state; // @[playground/src/cache/ICache.scala 327:53 328:15 92:94]
  wire [2:0] _GEN_1731 = io_cpu_tlb_hit ? 3'h0 : state; // @[playground/src/cache/ICache.scala 343:30 344:17 92:94]
  wire  _GEN_1732 = io_cpu_tlb_page_fault | page_fault; // @[playground/src/cache/ICache.scala 218:32 337:41 338:32]
  wire [2:0] _GEN_1733 = io_cpu_tlb_page_fault ? 3'h3 : _GEN_1731; // @[playground/src/cache/ICache.scala 337:41 339:32]
  wire [31:0] _GEN_1734 = io_cpu_tlb_page_fault ? 32'h13 : rdata_in_wait_0_inst; // @[playground/src/cache/ICache.scala 149:30 337:41 340:32]
  wire  _GEN_1735 = io_cpu_tlb_page_fault | rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 149:30 337:41 341:32]
  wire [2:0] _GEN_1742 = 3'h5 == state ? _GEN_1733 : state; // @[playground/src/cache/ICache.scala 233:17 92:94]
  wire [31:0] _GEN_1743 = 3'h5 == state ? _GEN_1734 : rdata_in_wait_0_inst; // @[playground/src/cache/ICache.scala 233:17 149:30]
  wire  _GEN_1744 = 3'h5 == state ? _GEN_1735 : rdata_in_wait_0_valid; // @[playground/src/cache/ICache.scala 233:17 149:30]
  wire  _GEN_1745 = 3'h5 == state ? _GEN_1732 : page_fault; // @[playground/src/cache/ICache.scala 233:17 218:32]
  wire [2:0] _GEN_1746 = 3'h4 == state ? _GEN_1730 : _GEN_1742; // @[playground/src/cache/ICache.scala 233:17]
  wire [31:0] _GEN_1748 = 3'h4 == state ? rdata_in_wait_0_inst : _GEN_1743; // @[playground/src/cache/ICache.scala 233:17 149:30]
  wire  _GEN_1749 = 3'h4 == state ? rdata_in_wait_0_valid : _GEN_1744; // @[playground/src/cache/ICache.scala 233:17 149:30]
  wire  _GEN_1750 = 3'h4 == state ? page_fault : _GEN_1745; // @[playground/src/cache/ICache.scala 233:17 218:32]
  wire  _GEN_1751 = 3'h3 == state ? _GEN_1724 : access_fault; // @[playground/src/cache/ICache.scala 233:17]
  wire  _GEN_1752 = 3'h3 == state ? _GEN_1725 : _GEN_1750; // @[playground/src/cache/ICache.scala 233:17]
  wire  _GEN_1753 = 3'h3 == state ? _GEN_1726 : addr_misaligned; // @[playground/src/cache/ICache.scala 233:17 219:32]
  wire [2:0] _GEN_1754 = 3'h3 == state ? _GEN_1727 : _GEN_1746; // @[playground/src/cache/ICache.scala 233:17]
  wire  _GEN_1755 = 3'h3 == state ? _GEN_1728 : _GEN_1749; // @[playground/src/cache/ICache.scala 233:17]
  wire  _GEN_1756 = 3'h3 == state ? _GEN_1729 : rdata_in_wait_1_valid; // @[playground/src/cache/ICache.scala 233:17 149:30]
  wire [31:0] _GEN_1757 = 3'h3 == state ? rdata_in_wait_0_inst : _GEN_1748; // @[playground/src/cache/ICache.scala 233:17 149:30]
  wire [2:0] _GEN_1778 = 3'h2 == state ? _GEN_1723 : _GEN_1754; // @[playground/src/cache/ICache.scala 233:17]
  SimpleDualPortRam bank_0_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_0_0_clock),
    .reset(bank_0_0_reset),
    .io_raddr(bank_0_0_io_raddr),
    .io_rdata(bank_0_0_io_rdata),
    .io_waddr(bank_0_0_io_waddr),
    .io_wen(bank_0_0_io_wen),
    .io_wstrb(bank_0_0_io_wstrb),
    .io_wdata(bank_0_0_io_wdata)
  );
  SimpleDualPortRam bank_1_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_1_0_clock),
    .reset(bank_1_0_reset),
    .io_raddr(bank_1_0_io_raddr),
    .io_rdata(bank_1_0_io_rdata),
    .io_waddr(bank_1_0_io_waddr),
    .io_wen(bank_1_0_io_wen),
    .io_wstrb(bank_1_0_io_wstrb),
    .io_wdata(bank_1_0_io_wdata)
  );
  SimpleDualPortRam bank_2_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_2_0_clock),
    .reset(bank_2_0_reset),
    .io_raddr(bank_2_0_io_raddr),
    .io_rdata(bank_2_0_io_rdata),
    .io_waddr(bank_2_0_io_waddr),
    .io_wen(bank_2_0_io_wen),
    .io_wstrb(bank_2_0_io_wstrb),
    .io_wdata(bank_2_0_io_wdata)
  );
  SimpleDualPortRam bank_3_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_3_0_clock),
    .reset(bank_3_0_reset),
    .io_raddr(bank_3_0_io_raddr),
    .io_rdata(bank_3_0_io_rdata),
    .io_waddr(bank_3_0_io_waddr),
    .io_wen(bank_3_0_io_wen),
    .io_wstrb(bank_3_0_io_wstrb),
    .io_wdata(bank_3_0_io_wdata)
  );
  SimpleDualPortRam bank_4_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_4_0_clock),
    .reset(bank_4_0_reset),
    .io_raddr(bank_4_0_io_raddr),
    .io_rdata(bank_4_0_io_rdata),
    .io_waddr(bank_4_0_io_waddr),
    .io_wen(bank_4_0_io_wen),
    .io_wstrb(bank_4_0_io_wstrb),
    .io_wdata(bank_4_0_io_wdata)
  );
  SimpleDualPortRam bank_5_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_5_0_clock),
    .reset(bank_5_0_reset),
    .io_raddr(bank_5_0_io_raddr),
    .io_rdata(bank_5_0_io_rdata),
    .io_waddr(bank_5_0_io_waddr),
    .io_wen(bank_5_0_io_wen),
    .io_wstrb(bank_5_0_io_wstrb),
    .io_wdata(bank_5_0_io_wdata)
  );
  SimpleDualPortRam bank_6_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_6_0_clock),
    .reset(bank_6_0_reset),
    .io_raddr(bank_6_0_io_raddr),
    .io_rdata(bank_6_0_io_rdata),
    .io_waddr(bank_6_0_io_waddr),
    .io_wen(bank_6_0_io_wen),
    .io_wstrb(bank_6_0_io_wstrb),
    .io_wdata(bank_6_0_io_wdata)
  );
  SimpleDualPortRam bank_7_0 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_7_0_clock),
    .reset(bank_7_0_reset),
    .io_raddr(bank_7_0_io_raddr),
    .io_rdata(bank_7_0_io_rdata),
    .io_waddr(bank_7_0_io_waddr),
    .io_wen(bank_7_0_io_wen),
    .io_wstrb(bank_7_0_io_wstrb),
    .io_wdata(bank_7_0_io_wdata)
  );
  SimpleDualPortRam bank_0_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_0_0_1_clock),
    .reset(bank_0_0_1_reset),
    .io_raddr(bank_0_0_1_io_raddr),
    .io_rdata(bank_0_0_1_io_rdata),
    .io_waddr(bank_0_0_1_io_waddr),
    .io_wen(bank_0_0_1_io_wen),
    .io_wstrb(bank_0_0_1_io_wstrb),
    .io_wdata(bank_0_0_1_io_wdata)
  );
  SimpleDualPortRam bank_1_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_1_0_1_clock),
    .reset(bank_1_0_1_reset),
    .io_raddr(bank_1_0_1_io_raddr),
    .io_rdata(bank_1_0_1_io_rdata),
    .io_waddr(bank_1_0_1_io_waddr),
    .io_wen(bank_1_0_1_io_wen),
    .io_wstrb(bank_1_0_1_io_wstrb),
    .io_wdata(bank_1_0_1_io_wdata)
  );
  SimpleDualPortRam bank_2_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_2_0_1_clock),
    .reset(bank_2_0_1_reset),
    .io_raddr(bank_2_0_1_io_raddr),
    .io_rdata(bank_2_0_1_io_rdata),
    .io_waddr(bank_2_0_1_io_waddr),
    .io_wen(bank_2_0_1_io_wen),
    .io_wstrb(bank_2_0_1_io_wstrb),
    .io_wdata(bank_2_0_1_io_wdata)
  );
  SimpleDualPortRam bank_3_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_3_0_1_clock),
    .reset(bank_3_0_1_reset),
    .io_raddr(bank_3_0_1_io_raddr),
    .io_rdata(bank_3_0_1_io_rdata),
    .io_waddr(bank_3_0_1_io_waddr),
    .io_wen(bank_3_0_1_io_wen),
    .io_wstrb(bank_3_0_1_io_wstrb),
    .io_wdata(bank_3_0_1_io_wdata)
  );
  SimpleDualPortRam bank_4_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_4_0_1_clock),
    .reset(bank_4_0_1_reset),
    .io_raddr(bank_4_0_1_io_raddr),
    .io_rdata(bank_4_0_1_io_rdata),
    .io_waddr(bank_4_0_1_io_waddr),
    .io_wen(bank_4_0_1_io_wen),
    .io_wstrb(bank_4_0_1_io_wstrb),
    .io_wdata(bank_4_0_1_io_wdata)
  );
  SimpleDualPortRam bank_5_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_5_0_1_clock),
    .reset(bank_5_0_1_reset),
    .io_raddr(bank_5_0_1_io_raddr),
    .io_rdata(bank_5_0_1_io_rdata),
    .io_waddr(bank_5_0_1_io_waddr),
    .io_wen(bank_5_0_1_io_wen),
    .io_wstrb(bank_5_0_1_io_wstrb),
    .io_wdata(bank_5_0_1_io_wdata)
  );
  SimpleDualPortRam bank_6_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_6_0_1_clock),
    .reset(bank_6_0_1_reset),
    .io_raddr(bank_6_0_1_io_raddr),
    .io_rdata(bank_6_0_1_io_rdata),
    .io_waddr(bank_6_0_1_io_waddr),
    .io_wen(bank_6_0_1_io_wen),
    .io_wstrb(bank_6_0_1_io_wstrb),
    .io_wdata(bank_6_0_1_io_wdata)
  );
  SimpleDualPortRam bank_7_0_1 ( // @[playground/src/cache/ICache.scala 168:17]
    .clock(bank_7_0_1_clock),
    .reset(bank_7_0_1_reset),
    .io_raddr(bank_7_0_1_io_raddr),
    .io_rdata(bank_7_0_1_io_rdata),
    .io_waddr(bank_7_0_1_io_waddr),
    .io_wen(bank_7_0_1_io_wen),
    .io_wstrb(bank_7_0_1_io_wstrb),
    .io_wdata(bank_7_0_1_io_wdata)
  );
  LUTRam tagBram ( // @[playground/src/cache/ICache.scala 192:25]
    .clock(tagBram_clock),
    .reset(tagBram_reset),
    .io_raddr(tagBram_io_raddr),
    .io_rdata(tagBram_io_rdata),
    .io_waddr(tagBram_io_waddr),
    .io_wdata(tagBram_io_wdata),
    .io_wen(tagBram_io_wen)
  );
  LUTRam tagBram_1 ( // @[playground/src/cache/ICache.scala 192:25]
    .clock(tagBram_1_clock),
    .reset(tagBram_1_reset),
    .io_raddr(tagBram_1_io_raddr),
    .io_rdata(tagBram_1_io_rdata),
    .io_waddr(tagBram_1_io_waddr),
    .io_wdata(tagBram_1_io_wdata),
    .io_wen(tagBram_1_io_wen)
  );
  assign io_cpu_inst_0 = {{32'd0}, _io_cpu_inst_0_T_1}; // @[playground/src/cache/ICache.scala 187:26]
  assign io_cpu_inst_1 = {{32'd0}, _io_cpu_inst_1_T_1}; // @[playground/src/cache/ICache.scala 187:26]
  assign io_cpu_inst_valid_0 = _io_cpu_inst_valid_0_T_1 & io_cpu_req; // @[playground/src/cache/ICache.scala 186:90]
  assign io_cpu_inst_valid_1 = _io_cpu_inst_valid_1_T_1 & io_cpu_req; // @[playground/src/cache/ICache.scala 186:90]
  assign io_cpu_access_fault = access_fault; // @[playground/src/cache/ICache.scala 229:26]
  assign io_cpu_page_fault = page_fault; // @[playground/src/cache/ICache.scala 230:26]
  assign io_cpu_addr_misaligned = addr_misaligned; // @[playground/src/cache/ICache.scala 231:26]
  assign io_cpu_icache_stall = _use_next_addr_T ? ~cache_hit_available & io_cpu_req : state != 3'h3; // @[playground/src/cache/ICache.scala 201:29]
  assign io_cpu_tlb_en = io_cpu_req & (_use_next_addr_T | state == 3'h5); // @[playground/src/cache/ICache.scala 205:52]
  assign io_cpu_tlb_vaddr = io_cpu_addr_0; // @[playground/src/cache/ICache.scala 203:38]
  assign io_cpu_tlb_complete_single_request = io_cpu_complete_single_request; // @[playground/src/cache/ICache.scala 204:38]
  assign io_axi_ar_valid = arvalid; // @[playground/src/cache/ICache.scala 210:11]
  assign io_axi_ar_bits_addr = ar_addr; // @[playground/src/cache/ICache.scala 209:6]
  assign io_axi_ar_bits_len = ar_len; // @[playground/src/cache/ICache.scala 209:6]
  assign io_axi_ar_bits_size = ar_size; // @[playground/src/cache/ICache.scala 209:6]
  assign io_axi_r_ready = rready; // @[playground/src/cache/ICache.scala 215:10]
  assign bank_0_0_clock = clock;
  assign bank_0_0_reset = reset;
  assign bank_0_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_0_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_0_0_io_wen = replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_0_0_io_wstrb = replace_wstrb_0_0_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_0_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_1_0_clock = clock;
  assign bank_1_0_reset = reset;
  assign bank_1_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_1_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_1_0_io_wen = replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_1_0_io_wstrb = replace_wstrb_0_1_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_1_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_2_0_clock = clock;
  assign bank_2_0_reset = reset;
  assign bank_2_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_2_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_2_0_io_wen = replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_2_0_io_wstrb = replace_wstrb_0_2_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_2_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_3_0_clock = clock;
  assign bank_3_0_reset = reset;
  assign bank_3_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_3_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_3_0_io_wen = replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_3_0_io_wstrb = replace_wstrb_0_3_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_3_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_4_0_clock = clock;
  assign bank_4_0_reset = reset;
  assign bank_4_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_4_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_4_0_io_wen = replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_4_0_io_wstrb = replace_wstrb_0_4_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_4_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_5_0_clock = clock;
  assign bank_5_0_reset = reset;
  assign bank_5_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_5_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_5_0_io_wen = replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_5_0_io_wstrb = replace_wstrb_0_5_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_5_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_6_0_clock = clock;
  assign bank_6_0_reset = reset;
  assign bank_6_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_6_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_6_0_io_wen = replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_6_0_io_wstrb = replace_wstrb_0_6_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_6_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_7_0_clock = clock;
  assign bank_7_0_reset = reset;
  assign bank_7_0_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_7_0_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_7_0_io_wen = replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_7_0_io_wstrb = replace_wstrb_0_7_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_7_0_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_0_0_1_clock = clock;
  assign bank_0_0_1_reset = reset;
  assign bank_0_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_0_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_0_0_1_io_wen = replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_0_0_1_io_wstrb = replace_wstrb_1_0_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_0_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_1_0_1_clock = clock;
  assign bank_1_0_1_reset = reset;
  assign bank_1_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_1_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_1_0_1_io_wen = replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_1_0_1_io_wstrb = replace_wstrb_1_1_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_1_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_2_0_1_clock = clock;
  assign bank_2_0_1_reset = reset;
  assign bank_2_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_2_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_2_0_1_io_wen = replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_2_0_1_io_wstrb = replace_wstrb_1_2_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_2_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_3_0_1_clock = clock;
  assign bank_3_0_1_reset = reset;
  assign bank_3_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_3_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_3_0_1_io_wen = replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_3_0_1_io_wstrb = replace_wstrb_1_3_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_3_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_4_0_1_clock = clock;
  assign bank_4_0_1_reset = reset;
  assign bank_4_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_4_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_4_0_1_io_wen = replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_4_0_1_io_wstrb = replace_wstrb_1_4_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_4_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_5_0_1_clock = clock;
  assign bank_5_0_1_reset = reset;
  assign bank_5_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_5_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_5_0_1_io_wen = replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_5_0_1_io_wstrb = replace_wstrb_1_5_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_5_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_6_0_1_clock = clock;
  assign bank_6_0_1_reset = reset;
  assign bank_6_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_6_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_6_0_1_io_wen = replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_6_0_1_io_wstrb = replace_wstrb_1_6_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_6_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign bank_7_0_1_clock = clock;
  assign bank_7_0_1_reset = reset;
  assign bank_7_0_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 102:47]
  assign bank_7_0_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign bank_7_0_1_io_wen = replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 177:29]
  assign bank_7_0_1_io_wstrb = replace_wstrb_1_7_0; // @[playground/src/cache/ICache.scala 180:29]
  assign bank_7_0_1_io_wdata = io_axi_r_bits_data; // @[playground/src/cache/ICache.scala 179:29]
  assign tagBram_clock = clock;
  assign tagBram_reset = reset;
  assign tagBram_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 105:45]
  assign tagBram_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign tagBram_io_wdata = tag_wdata; // @[playground/src/cache/ICache.scala 198:22]
  assign tagBram_io_wen = tag_wstrb_0; // @[playground/src/cache/ICache.scala 196:22]
  assign tagBram_1_clock = clock;
  assign tagBram_1_reset = reset;
  assign tagBram_1_io_raddr = _GEN_1[11:6]; // @[playground/src/cache/ICache.scala 105:45]
  assign tagBram_1_io_waddr = io_cpu_addr_0[11:6]; // @[playground/src/cache/ICache.scala 112:37]
  assign tagBram_1_io_wdata = tag_wdata; // @[playground/src/cache/ICache.scala 198:22]
  assign tagBram_1_io_wen = tag_wstrb_1; // @[playground/src/cache/ICache.scala 196:22]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/cache/ICache.scala 92:94]
      state <= 3'h0; // @[playground/src/cache/ICache.scala 92:94]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      state <= 3'h4; // @[playground/src/cache/ICache.scala 354:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        state <= _GEN_1159;
      end
    end else if (3'h1 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      state <= _GEN_1613;
    end else begin
      state <= _GEN_1778;
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_0 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_0 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_0 <= _GEN_1185;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_1 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_1 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_1 <= _GEN_1186;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_2 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_2 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_2 <= _GEN_1187;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_3 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_3 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_3 <= _GEN_1188;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_4 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_4 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_4 <= _GEN_1189;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_5 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_5 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_5 <= _GEN_1190;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_6 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_6 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_6 <= _GEN_1191;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_7 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_7 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_7 <= _GEN_1192;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_8 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_8 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_8 <= _GEN_1193;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_9 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_9 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_9 <= _GEN_1194;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_10 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_10 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_10 <= _GEN_1195;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_11 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_11 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_11 <= _GEN_1196;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_12 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_12 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_12 <= _GEN_1197;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_13 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_13 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_13 <= _GEN_1198;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_14 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_14 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_14 <= _GEN_1199;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_15 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_15 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_15 <= _GEN_1200;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_16 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_16 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_16 <= _GEN_1201;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_17 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_17 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_17 <= _GEN_1202;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_18 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_18 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_18 <= _GEN_1203;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_19 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_19 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_19 <= _GEN_1204;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_20 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_20 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_20 <= _GEN_1205;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_21 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_21 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_21 <= _GEN_1206;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_22 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_22 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_22 <= _GEN_1207;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_23 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_23 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_23 <= _GEN_1208;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_24 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_24 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_24 <= _GEN_1209;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_25 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_25 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_25 <= _GEN_1210;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_26 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_26 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_26 <= _GEN_1211;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_27 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_27 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_27 <= _GEN_1212;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_28 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_28 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_28 <= _GEN_1213;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_29 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_29 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_29 <= _GEN_1214;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_30 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_30 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_30 <= _GEN_1215;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_31 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_31 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_31 <= _GEN_1216;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_32 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_32 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_32 <= _GEN_1217;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_33 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_33 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_33 <= _GEN_1218;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_34 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_34 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_34 <= _GEN_1219;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_35 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_35 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_35 <= _GEN_1220;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_36 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_36 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_36 <= _GEN_1221;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_37 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_37 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_37 <= _GEN_1222;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_38 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_38 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_38 <= _GEN_1223;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_39 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_39 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_39 <= _GEN_1224;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_40 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_40 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_40 <= _GEN_1225;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_41 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_41 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_41 <= _GEN_1226;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_42 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_42 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_42 <= _GEN_1227;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_43 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_43 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_43 <= _GEN_1228;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_44 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_44 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_44 <= _GEN_1229;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_45 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_45 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_45 <= _GEN_1230;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_46 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_46 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_46 <= _GEN_1231;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_47 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_47 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_47 <= _GEN_1232;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_48 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_48 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_48 <= _GEN_1233;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_49 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_49 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_49 <= _GEN_1234;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_50 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_50 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_50 <= _GEN_1235;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_51 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_51 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_51 <= _GEN_1236;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_52 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_52 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_52 <= _GEN_1237;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_53 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_53 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_53 <= _GEN_1238;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_54 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_54 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_54 <= _GEN_1239;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_55 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_55 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_55 <= _GEN_1240;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_56 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_56 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_56 <= _GEN_1241;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_57 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_57 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_57 <= _GEN_1242;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_58 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_58 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_58 <= _GEN_1243;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_59 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_59 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_59 <= _GEN_1244;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_60 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_60 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_60 <= _GEN_1245;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_61 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_61 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_61 <= _GEN_1246;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_62 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_62 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_62 <= _GEN_1247;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_0_63 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_0_63 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_0_63 <= _GEN_1248;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_0 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_0 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_0 <= _GEN_1249;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_1 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_1 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_1 <= _GEN_1250;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_2 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_2 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_2 <= _GEN_1251;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_3 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_3 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_3 <= _GEN_1252;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_4 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_4 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_4 <= _GEN_1253;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_5 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_5 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_5 <= _GEN_1254;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_6 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_6 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_6 <= _GEN_1255;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_7 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_7 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_7 <= _GEN_1256;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_8 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_8 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_8 <= _GEN_1257;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_9 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_9 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_9 <= _GEN_1258;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_10 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_10 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_10 <= _GEN_1259;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_11 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_11 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_11 <= _GEN_1260;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_12 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_12 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_12 <= _GEN_1261;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_13 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_13 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_13 <= _GEN_1262;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_14 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_14 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_14 <= _GEN_1263;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_15 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_15 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_15 <= _GEN_1264;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_16 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_16 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_16 <= _GEN_1265;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_17 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_17 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_17 <= _GEN_1266;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_18 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_18 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_18 <= _GEN_1267;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_19 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_19 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_19 <= _GEN_1268;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_20 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_20 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_20 <= _GEN_1269;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_21 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_21 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_21 <= _GEN_1270;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_22 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_22 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_22 <= _GEN_1271;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_23 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_23 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_23 <= _GEN_1272;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_24 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_24 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_24 <= _GEN_1273;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_25 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_25 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_25 <= _GEN_1274;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_26 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_26 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_26 <= _GEN_1275;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_27 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_27 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_27 <= _GEN_1276;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_28 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_28 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_28 <= _GEN_1277;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_29 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_29 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_29 <= _GEN_1278;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_30 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_30 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_30 <= _GEN_1279;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_31 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_31 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_31 <= _GEN_1280;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_32 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_32 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_32 <= _GEN_1281;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_33 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_33 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_33 <= _GEN_1282;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_34 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_34 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_34 <= _GEN_1283;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_35 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_35 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_35 <= _GEN_1284;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_36 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_36 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_36 <= _GEN_1285;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_37 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_37 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_37 <= _GEN_1286;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_38 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_38 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_38 <= _GEN_1287;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_39 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_39 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_39 <= _GEN_1288;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_40 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_40 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_40 <= _GEN_1289;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_41 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_41 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_41 <= _GEN_1290;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_42 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_42 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_42 <= _GEN_1291;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_43 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_43 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_43 <= _GEN_1292;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_44 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_44 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_44 <= _GEN_1293;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_45 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_45 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_45 <= _GEN_1294;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_46 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_46 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_46 <= _GEN_1295;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_47 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_47 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_47 <= _GEN_1296;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_48 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_48 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_48 <= _GEN_1297;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_49 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_49 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_49 <= _GEN_1298;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_50 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_50 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_50 <= _GEN_1299;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_51 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_51 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_51 <= _GEN_1300;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_52 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_52 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_52 <= _GEN_1301;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_53 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_53 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_53 <= _GEN_1302;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_54 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_54 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_54 <= _GEN_1303;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_55 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_55 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_55 <= _GEN_1304;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_56 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_56 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_56 <= _GEN_1305;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_57 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_57 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_57 <= _GEN_1306;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_58 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_58 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_58 <= _GEN_1307;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_59 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_59 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_59 <= _GEN_1308;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_60 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_60 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_60 <= _GEN_1309;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_61 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_61 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_61 <= _GEN_1310;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_62 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_62 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_62 <= _GEN_1311;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 95:22]
      valid_1_63 <= 1'h0; // @[playground/src/cache/ICache.scala 95:22]
    end else if (io_cpu_fence_i) begin // @[playground/src/cache/ICache.scala 352:24]
      valid_1_63 <= 1'h0; // @[playground/src/cache/ICache.scala 353:11]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        valid_1_63 <= _GEN_1312;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 104:26]
      tag_0 <= 20'h0; // @[playground/src/cache/ICache.scala 104:26]
    end else begin
      tag_0 <= tagBram_io_rdata; // @[playground/src/cache/ICache.scala 194:22]
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 104:26]
      tag_1 <= 20'h0; // @[playground/src/cache/ICache.scala 104:26]
    end else begin
      tag_1 <= tagBram_1_io_rdata; // @[playground/src/cache/ICache.scala 194:22]
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 106:26]
      tag_wstrb_0 <= 1'h0; // @[playground/src/cache/ICache.scala 106:26]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          tag_wstrb_0 <= _GEN_959;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        tag_wstrb_0 <= _GEN_1721;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 106:26]
      tag_wstrb_1 <= 1'h0; // @[playground/src/cache/ICache.scala 106:26]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          tag_wstrb_1 <= _GEN_960;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        tag_wstrb_1 <= _GEN_1722;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 107:26]
      tag_wdata <= 20'h0; // @[playground/src/cache/ICache.scala 107:26]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          tag_wdata <= _GEN_961;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_0 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_0 <= _GEN_1090;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_1 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_1 <= _GEN_1091;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_2 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_2 <= _GEN_1092;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_3 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_3 <= _GEN_1093;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_4 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_4 <= _GEN_1094;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_5 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_5 <= _GEN_1095;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_6 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_6 <= _GEN_1096;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_7 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_7 <= _GEN_1097;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_8 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_8 <= _GEN_1098;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_9 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_9 <= _GEN_1099;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_10 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_10 <= _GEN_1100;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_11 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_11 <= _GEN_1101;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_12 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_12 <= _GEN_1102;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_13 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_13 <= _GEN_1103;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_14 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_14 <= _GEN_1104;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_15 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_15 <= _GEN_1105;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_16 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_16 <= _GEN_1106;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_17 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_17 <= _GEN_1107;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_18 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_18 <= _GEN_1108;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_19 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_19 <= _GEN_1109;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_20 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_20 <= _GEN_1110;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_21 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_21 <= _GEN_1111;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_22 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_22 <= _GEN_1112;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_23 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_23 <= _GEN_1113;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_24 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_24 <= _GEN_1114;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_25 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_25 <= _GEN_1115;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_26 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_26 <= _GEN_1116;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_27 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_27 <= _GEN_1117;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_28 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_28 <= _GEN_1118;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_29 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_29 <= _GEN_1119;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_30 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_30 <= _GEN_1120;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_31 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_31 <= _GEN_1121;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_32 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_32 <= _GEN_1122;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_33 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_33 <= _GEN_1123;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_34 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_34 <= _GEN_1124;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_35 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_35 <= _GEN_1125;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_36 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_36 <= _GEN_1126;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_37 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_37 <= _GEN_1127;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_38 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_38 <= _GEN_1128;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_39 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_39 <= _GEN_1129;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_40 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_40 <= _GEN_1130;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_41 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_41 <= _GEN_1131;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_42 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_42 <= _GEN_1132;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_43 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_43 <= _GEN_1133;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_44 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_44 <= _GEN_1134;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_45 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_45 <= _GEN_1135;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_46 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_46 <= _GEN_1136;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_47 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_47 <= _GEN_1137;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_48 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_48 <= _GEN_1138;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_49 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_49 <= _GEN_1139;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_50 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_50 <= _GEN_1140;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_51 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_51 <= _GEN_1141;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_52 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_52 <= _GEN_1142;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_53 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_53 <= _GEN_1143;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_54 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_54 <= _GEN_1144;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_55 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_55 <= _GEN_1145;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_56 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_56 <= _GEN_1146;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_57 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_57 <= _GEN_1147;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_58 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_58 <= _GEN_1148;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_59 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_59 <= _GEN_1149;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_60 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_60 <= _GEN_1150;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_61 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_61 <= _GEN_1151;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_62 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_62 <= _GEN_1152;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 110:20]
      lru_63 <= 1'h0; // @[playground/src/cache/ICache.scala 110:20]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          lru_63 <= _GEN_1153;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_0_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_0_0 <= _GEN_943;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_0_0 <= _GEN_1705;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_1_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_1_0 <= _GEN_945;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_1_0 <= _GEN_1707;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_2_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_2_0 <= _GEN_947;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_2_0 <= _GEN_1709;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_3_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_3_0 <= _GEN_949;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_3_0 <= _GEN_1711;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_4_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_4_0 <= _GEN_951;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_4_0 <= _GEN_1713;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_5_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_5_0 <= _GEN_953;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_5_0 <= _GEN_1715;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_6_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_6_0 <= _GEN_955;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_6_0 <= _GEN_1717;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_0_7_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_0_7_0 <= _GEN_957;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_0_7_0 <= _GEN_1719;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_0_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_0_0 <= _GEN_944;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_0_0 <= _GEN_1706;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_1_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_1_0 <= _GEN_946;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_1_0 <= _GEN_1708;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_2_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_2_0 <= _GEN_948;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_2_0 <= _GEN_1710;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_3_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_3_0 <= _GEN_950;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_3_0 <= _GEN_1712;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_4_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_4_0 <= _GEN_952;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_4_0 <= _GEN_1714;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_5_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_5_0 <= _GEN_954;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_5_0 <= _GEN_1716;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_6_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_6_0 <= _GEN_956;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_6_0 <= _GEN_1718;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 117:30]
      replace_wstrb_1_7_0 <= 1'h0; // @[playground/src/cache/ICache.scala 117:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          replace_wstrb_1_7_0 <= _GEN_958;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        replace_wstrb_1_7_0 <= _GEN_1720;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 149:30]
      rdata_in_wait_0_inst <= 32'h0; // @[playground/src/cache/ICache.scala 149:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (addr_err) begin // @[playground/src/cache/ICache.scala 239:24]
          rdata_in_wait_0_inst <= 32'h13; // @[playground/src/cache/ICache.scala 246:34]
        end
      end
    end else if (3'h1 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (!(io_axi_ar_valid)) begin // @[playground/src/cache/ICache.scala 280:29]
        rdata_in_wait_0_inst <= _GEN_1603;
      end
    end else if (!(3'h2 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      rdata_in_wait_0_inst <= _GEN_1757;
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 149:30]
      rdata_in_wait_0_valid <= 1'h0; // @[playground/src/cache/ICache.scala 149:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        rdata_in_wait_0_valid <= _GEN_1161;
      end
    end else if (3'h1 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (!(io_axi_ar_valid)) begin // @[playground/src/cache/ICache.scala 280:29]
        rdata_in_wait_0_valid <= _GEN_1604;
      end
    end else if (!(3'h2 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      rdata_in_wait_0_valid <= _GEN_1755;
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 149:30]
      rdata_in_wait_1_inst <= 32'h0; // @[playground/src/cache/ICache.scala 149:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          rdata_in_wait_1_inst <= _GEN_1154;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 149:30]
      rdata_in_wait_1_valid <= 1'h0; // @[playground/src/cache/ICache.scala 149:30]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          rdata_in_wait_1_valid <= _GEN_1156;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (!(3'h2 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
        rdata_in_wait_1_valid <= _GEN_1756;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 207:24]
      ar_addr <= 32'h0; // @[playground/src/cache/ICache.scala 207:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          ar_addr <= _GEN_939;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 207:24]
      ar_len <= 8'h0; // @[playground/src/cache/ICache.scala 207:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          ar_len <= _GEN_940;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 207:24]
      ar_size <= 3'h0; // @[playground/src/cache/ICache.scala 207:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          ar_size <= _GEN_941;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 208:24]
      arvalid <= 1'h0; // @[playground/src/cache/ICache.scala 208:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (io_cpu_req) begin // @[playground/src/cache/ICache.scala 238:24]
        if (!(addr_err)) begin // @[playground/src/cache/ICache.scala 239:24]
          arvalid <= _GEN_942;
        end
      end
    end else if (3'h1 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      arvalid <= _GEN_1608;
    end else if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      arvalid <= _GEN_1608;
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 213:23]
      rready <= 1'h0; // @[playground/src/cache/ICache.scala 213:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (3'h1 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        if (io_axi_ar_valid) begin // @[playground/src/cache/ICache.scala 280:29]
          rready <= _GEN_1602;
        end else begin
          rready <= _GEN_1605;
        end
      end else if (3'h2 == state) begin // @[playground/src/cache/ICache.scala 233:17]
        rready <= _GEN_1704;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 217:32]
      access_fault <= 1'h0; // @[playground/src/cache/ICache.scala 217:32]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      access_fault <= _GEN_1380;
    end else if (3'h1 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      if (!(io_axi_ar_valid)) begin // @[playground/src/cache/ICache.scala 280:29]
        access_fault <= _GEN_1606;
      end
    end else if (!(3'h2 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      access_fault <= _GEN_1751;
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 218:32]
      page_fault <= 1'h0; // @[playground/src/cache/ICache.scala 218:32]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      page_fault <= 1'h0; // @[playground/src/cache/ICache.scala 236:23]
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (!(3'h2 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
        page_fault <= _GEN_1752;
      end
    end
    if (reset) begin // @[playground/src/cache/ICache.scala 219:32]
      addr_misaligned <= 1'h0; // @[playground/src/cache/ICache.scala 219:32]
    end else if (3'h0 == state) begin // @[playground/src/cache/ICache.scala 233:17]
      addr_misaligned <= _GEN_1379;
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
      if (!(3'h2 == state)) begin // @[playground/src/cache/ICache.scala 233:17]
        addr_misaligned <= _GEN_1753;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  valid_0_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_0_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_0_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_0_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_0_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_0_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_0_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_0_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_0_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_0_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_0_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_0_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_0_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_0_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_0_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_0_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_0_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_0_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_0_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_0_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_0_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_0_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_0_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_0_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_0_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_0_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_0_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_0_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_0_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_0_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_0_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_0_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_0_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_0_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_0_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_0_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_0_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_0_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_0_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_0_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_0_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_0_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_0_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_0_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_0_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_0_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_0_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_0_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_0_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_0_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_0_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_0_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_0_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_0_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_0_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_0_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_0_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_0_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_0_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_0_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_0_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_0_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_0_62 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_0_63 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_1_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_1_1 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_1_2 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_1_3 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_1_4 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_1_5 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_1_6 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_1_7 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_1_8 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_1_9 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_1_10 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_1_11 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_1_12 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_1_13 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_1_14 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_1_15 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1_16 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_1_17 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_18 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_1_19 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_1_20 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_1_21 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_1_22 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_1_23 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_1_24 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_1_25 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_1_26 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_1_27 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_1_28 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_1_29 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_1_30 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_1_31 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_1_32 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_1_33 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_1_34 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_1_35 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_1_36 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_1_37 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_1_38 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_1_39 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_1_40 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_1_41 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_1_42 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_1_43 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_1_44 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_1_45 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_1_46 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_1_47 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_1_48 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_1_49 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_1_50 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_1_51 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_1_52 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_1_53 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_1_54 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_1_55 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_1_56 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_1_57 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_1_58 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_1_59 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_1_60 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_1_61 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_1_62 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_1_63 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  tag_0 = _RAND_129[19:0];
  _RAND_130 = {1{`RANDOM}};
  tag_1 = _RAND_130[19:0];
  _RAND_131 = {1{`RANDOM}};
  tag_wstrb_0 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  tag_wstrb_1 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  tag_wdata = _RAND_133[19:0];
  _RAND_134 = {1{`RANDOM}};
  lru_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  lru_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  lru_2 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  lru_3 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  lru_4 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  lru_5 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  lru_6 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  lru_7 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  lru_8 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  lru_9 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  lru_10 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  lru_11 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  lru_12 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  lru_13 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  lru_14 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  lru_15 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  lru_16 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  lru_17 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  lru_18 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  lru_19 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  lru_20 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  lru_21 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  lru_22 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  lru_23 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  lru_24 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  lru_25 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  lru_26 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  lru_27 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  lru_28 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  lru_29 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  lru_30 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  lru_31 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  lru_32 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  lru_33 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  lru_34 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  lru_35 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  lru_36 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  lru_37 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  lru_38 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  lru_39 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  lru_40 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  lru_41 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  lru_42 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  lru_43 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  lru_44 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  lru_45 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  lru_46 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  lru_47 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  lru_48 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  lru_49 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  lru_50 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  lru_51 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  lru_52 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  lru_53 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  lru_54 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  lru_55 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  lru_56 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  lru_57 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  lru_58 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  lru_59 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  lru_60 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  lru_61 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  lru_62 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  lru_63 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  replace_wstrb_0_0_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  replace_wstrb_0_1_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  replace_wstrb_0_2_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  replace_wstrb_0_3_0 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  replace_wstrb_0_4_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  replace_wstrb_0_5_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  replace_wstrb_0_6_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  replace_wstrb_0_7_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  replace_wstrb_1_0_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  replace_wstrb_1_1_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  replace_wstrb_1_2_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  replace_wstrb_1_3_0 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  replace_wstrb_1_4_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  replace_wstrb_1_5_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  replace_wstrb_1_6_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  replace_wstrb_1_7_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  rdata_in_wait_0_inst = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  rdata_in_wait_0_valid = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  rdata_in_wait_1_inst = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  rdata_in_wait_1_valid = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ar_addr = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  ar_len = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  ar_size = _RAND_220[2:0];
  _RAND_221 = {1{`RANDOM}};
  arvalid = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  rready = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  access_fault = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  page_fault = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  addr_misaligned = _RAND_225[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [63:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [7:0]  io_enq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [63:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [7:0]  io_deq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [2:0]  io_deq_bits_size // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [63:0] ram_addr [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [7:0] ram_strb [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_strb_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [7:0] ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_strb_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_strb_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_strb_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [2:0] ram_size [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [1:0] ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 278:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 279:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 280:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = enq_ptr_value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 304:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 303:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 287:16]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 291:16]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 294:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 295:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_strb[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enq_ptr_value = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  deq_ptr_value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleDualPortRam_16(
  input         clock,
  input         reset,
  input  [5:0]  io_raddr, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  output [63:0] io_rdata, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input  [5:0]  io_waddr, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input         io_wen, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input  [7:0]  io_wstrb, // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
  input  [63:0] io_wdata // @[playground/src/cache/memory/SimpleDualPortRam.scala 34:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] bank_0 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_0_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_0_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_0_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_0_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_0_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_0_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_0_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_0_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_0_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_1 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_1_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_1_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_1_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_1_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_1_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_1_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_1_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_1_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_1_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_2 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_2_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_2_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_2_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_2_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_2_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_2_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_2_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_2_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_2_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_3 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_3_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_3_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_3_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_3_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_3_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_3_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_3_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_3_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_3_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_4 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_4_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_4_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_4_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_4_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_4_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_4_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_4_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_4_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_4_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_5 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_5_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_5_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_5_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_5_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_5_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_5_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_5_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_5_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_5_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_6 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_6_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_6_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_6_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_6_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_6_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_6_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_6_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_6_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_6_io_rdata_MPORT_addr_pipe_0;
  reg [7:0] bank_7 [0:63]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_7_io_rdata_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_7_io_rdata_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_7_io_rdata_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [7:0] bank_7_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire [5:0] bank_7_MPORT_addr; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_7_MPORT_mask; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  wire  bank_7_MPORT_en; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  reg  bank_7_io_rdata_MPORT_en_pipe_0;
  reg [5:0] bank_7_io_rdata_MPORT_addr_pipe_0;
  wire  _T_2 = |io_wstrb | ~io_wen; // @[playground/src/cache/memory/SimpleDualPortRam.scala 69:20]
  wire [31:0] io_rdata_lo = {bank_3_io_rdata_MPORT_data,bank_2_io_rdata_MPORT_data,bank_1_io_rdata_MPORT_data,
    bank_0_io_rdata_MPORT_data}; // @[playground/src/cache/memory/SimpleDualPortRam.scala 75:49]
  wire [31:0] io_rdata_hi = {bank_7_io_rdata_MPORT_data,bank_6_io_rdata_MPORT_data,bank_5_io_rdata_MPORT_data,
    bank_4_io_rdata_MPORT_data}; // @[playground/src/cache/memory/SimpleDualPortRam.scala 75:49]
  assign bank_0_io_rdata_MPORT_en = bank_0_io_rdata_MPORT_en_pipe_0;
  assign bank_0_io_rdata_MPORT_addr = bank_0_io_rdata_MPORT_addr_pipe_0;
  assign bank_0_io_rdata_MPORT_data = bank_0[bank_0_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_0_MPORT_data = io_wdata[7:0];
  assign bank_0_MPORT_addr = io_waddr;
  assign bank_0_MPORT_mask = io_wstrb[0];
  assign bank_0_MPORT_en = io_wen;
  assign bank_1_io_rdata_MPORT_en = bank_1_io_rdata_MPORT_en_pipe_0;
  assign bank_1_io_rdata_MPORT_addr = bank_1_io_rdata_MPORT_addr_pipe_0;
  assign bank_1_io_rdata_MPORT_data = bank_1[bank_1_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_1_MPORT_data = io_wdata[15:8];
  assign bank_1_MPORT_addr = io_waddr;
  assign bank_1_MPORT_mask = io_wstrb[1];
  assign bank_1_MPORT_en = io_wen;
  assign bank_2_io_rdata_MPORT_en = bank_2_io_rdata_MPORT_en_pipe_0;
  assign bank_2_io_rdata_MPORT_addr = bank_2_io_rdata_MPORT_addr_pipe_0;
  assign bank_2_io_rdata_MPORT_data = bank_2[bank_2_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_2_MPORT_data = io_wdata[23:16];
  assign bank_2_MPORT_addr = io_waddr;
  assign bank_2_MPORT_mask = io_wstrb[2];
  assign bank_2_MPORT_en = io_wen;
  assign bank_3_io_rdata_MPORT_en = bank_3_io_rdata_MPORT_en_pipe_0;
  assign bank_3_io_rdata_MPORT_addr = bank_3_io_rdata_MPORT_addr_pipe_0;
  assign bank_3_io_rdata_MPORT_data = bank_3[bank_3_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_3_MPORT_data = io_wdata[31:24];
  assign bank_3_MPORT_addr = io_waddr;
  assign bank_3_MPORT_mask = io_wstrb[3];
  assign bank_3_MPORT_en = io_wen;
  assign bank_4_io_rdata_MPORT_en = bank_4_io_rdata_MPORT_en_pipe_0;
  assign bank_4_io_rdata_MPORT_addr = bank_4_io_rdata_MPORT_addr_pipe_0;
  assign bank_4_io_rdata_MPORT_data = bank_4[bank_4_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_4_MPORT_data = io_wdata[39:32];
  assign bank_4_MPORT_addr = io_waddr;
  assign bank_4_MPORT_mask = io_wstrb[4];
  assign bank_4_MPORT_en = io_wen;
  assign bank_5_io_rdata_MPORT_en = bank_5_io_rdata_MPORT_en_pipe_0;
  assign bank_5_io_rdata_MPORT_addr = bank_5_io_rdata_MPORT_addr_pipe_0;
  assign bank_5_io_rdata_MPORT_data = bank_5[bank_5_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_5_MPORT_data = io_wdata[47:40];
  assign bank_5_MPORT_addr = io_waddr;
  assign bank_5_MPORT_mask = io_wstrb[5];
  assign bank_5_MPORT_en = io_wen;
  assign bank_6_io_rdata_MPORT_en = bank_6_io_rdata_MPORT_en_pipe_0;
  assign bank_6_io_rdata_MPORT_addr = bank_6_io_rdata_MPORT_addr_pipe_0;
  assign bank_6_io_rdata_MPORT_data = bank_6[bank_6_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_6_MPORT_data = io_wdata[55:48];
  assign bank_6_MPORT_addr = io_waddr;
  assign bank_6_MPORT_mask = io_wstrb[6];
  assign bank_6_MPORT_en = io_wen;
  assign bank_7_io_rdata_MPORT_en = bank_7_io_rdata_MPORT_en_pipe_0;
  assign bank_7_io_rdata_MPORT_addr = bank_7_io_rdata_MPORT_addr_pipe_0;
  assign bank_7_io_rdata_MPORT_data = bank_7[bank_7_io_rdata_MPORT_addr]; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
  assign bank_7_MPORT_data = io_wdata[63:56];
  assign bank_7_MPORT_addr = io_waddr;
  assign bank_7_MPORT_mask = io_wstrb[7];
  assign bank_7_MPORT_en = io_wen;
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[playground/src/cache/memory/SimpleDualPortRam.scala 75:49]
  always @(posedge clock) begin
    if (bank_0_MPORT_en & bank_0_MPORT_mask) begin
      bank_0[bank_0_MPORT_addr] <= bank_0_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_0_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_0_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_1_MPORT_en & bank_1_MPORT_mask) begin
      bank_1[bank_1_MPORT_addr] <= bank_1_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_1_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_1_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_2_MPORT_en & bank_2_MPORT_mask) begin
      bank_2[bank_2_MPORT_addr] <= bank_2_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_2_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_2_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_3_MPORT_en & bank_3_MPORT_mask) begin
      bank_3[bank_3_MPORT_addr] <= bank_3_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_3_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_3_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_4_MPORT_en & bank_4_MPORT_mask) begin
      bank_4[bank_4_MPORT_addr] <= bank_4_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_4_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_4_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_5_MPORT_en & bank_5_MPORT_mask) begin
      bank_5[bank_5_MPORT_addr] <= bank_5_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_5_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_5_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_6_MPORT_en & bank_6_MPORT_mask) begin
      bank_6[bank_6_MPORT_addr] <= bank_6_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_6_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_6_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    if (bank_7_MPORT_en & bank_7_MPORT_mask) begin
      bank_7[bank_7_MPORT_addr] <= bank_7_MPORT_data; // @[playground/src/cache/memory/SimpleDualPortRam.scala 73:29]
    end
    bank_7_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      bank_7_io_rdata_MPORT_addr_pipe_0 <= io_raddr;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed: when write port enable is high, write vector cannot be all 0\n    at SimpleDualPortRam.scala:68 assert(\n"
            ); // @[playground/src/cache/memory/SimpleDualPortRam.scala 68:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~_T_2) begin
          $fatal; // @[playground/src/cache/memory/SimpleDualPortRam.scala 68:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_3[initvar] = _RAND_9[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_4[initvar] = _RAND_12[7:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_5[initvar] = _RAND_15[7:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_6[initvar] = _RAND_18[7:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bank_7[initvar] = _RAND_21[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bank_0_io_rdata_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_4 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  bank_1_io_rdata_MPORT_addr_pipe_0 = _RAND_5[5:0];
  _RAND_7 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  bank_2_io_rdata_MPORT_addr_pipe_0 = _RAND_8[5:0];
  _RAND_10 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bank_3_io_rdata_MPORT_addr_pipe_0 = _RAND_11[5:0];
  _RAND_13 = {1{`RANDOM}};
  bank_4_io_rdata_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bank_4_io_rdata_MPORT_addr_pipe_0 = _RAND_14[5:0];
  _RAND_16 = {1{`RANDOM}};
  bank_5_io_rdata_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  bank_5_io_rdata_MPORT_addr_pipe_0 = _RAND_17[5:0];
  _RAND_19 = {1{`RANDOM}};
  bank_6_io_rdata_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  bank_6_io_rdata_MPORT_addr_pipe_0 = _RAND_20[5:0];
  _RAND_22 = {1{`RANDOM}};
  bank_7_io_rdata_MPORT_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  bank_7_io_rdata_MPORT_addr_pipe_0 = _RAND_23[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input         clock,
  input         reset,
  input  [63:0] io_cpu_exe_addr, // @[playground/src/cache/DCache.scala 83:14]
  input  [63:0] io_cpu_addr, // @[playground/src/cache/DCache.scala 83:14]
  input  [7:0]  io_cpu_rlen, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_en, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_wen, // @[playground/src/cache/DCache.scala 83:14]
  input  [63:0] io_cpu_wdata, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_complete_single_request, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_fence_i, // @[playground/src/cache/DCache.scala 83:14]
  input  [7:0]  io_cpu_wstrb, // @[playground/src/cache/DCache.scala 83:14]
  output [63:0] io_cpu_rdata, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_access_fault, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_page_fault, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_dcache_ready, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_en, // @[playground/src/cache/DCache.scala 83:14]
  output [63:0] io_cpu_tlb_vaddr, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_complete_single_request, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_tlb_uncached, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_tlb_hit, // @[playground/src/cache/DCache.scala 83:14]
  input  [19:0] io_cpu_tlb_ptag, // @[playground/src/cache/DCache.scala 83:14]
  input  [31:0] io_cpu_tlb_paddr, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_tlb_page_fault, // @[playground/src/cache/DCache.scala 83:14]
  output [1:0]  io_cpu_tlb_access_type, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_vpn_ready, // @[playground/src/cache/DCache.scala 83:14]
  input         io_cpu_tlb_ptw_vpn_valid, // @[playground/src/cache/DCache.scala 83:14]
  input  [26:0] io_cpu_tlb_ptw_vpn_bits, // @[playground/src/cache/DCache.scala 83:14]
  input  [1:0]  io_cpu_tlb_ptw_access_type, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_valid, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_access_fault, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_page_fault, // @[playground/src/cache/DCache.scala 83:14]
  output [19:0] io_cpu_tlb_ptw_pte_bits_entry_ppn, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_d, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_g, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_u, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_x, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_w, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_r, // @[playground/src/cache/DCache.scala 83:14]
  output        io_cpu_tlb_ptw_pte_bits_entry_flag_v, // @[playground/src/cache/DCache.scala 83:14]
  output [17:0] io_cpu_tlb_ptw_pte_bits_rmask, // @[playground/src/cache/DCache.scala 83:14]
  input  [63:0] io_cpu_tlb_csr_satp, // @[playground/src/cache/DCache.scala 83:14]
  input  [63:0] io_cpu_tlb_csr_mstatus, // @[playground/src/cache/DCache.scala 83:14]
  input  [1:0]  io_cpu_tlb_csr_imode, // @[playground/src/cache/DCache.scala 83:14]
  input  [1:0]  io_cpu_tlb_csr_dmode, // @[playground/src/cache/DCache.scala 83:14]
  input         io_axi_ar_ready, // @[playground/src/cache/DCache.scala 83:14]
  output        io_axi_ar_valid, // @[playground/src/cache/DCache.scala 83:14]
  output [31:0] io_axi_ar_bits_addr, // @[playground/src/cache/DCache.scala 83:14]
  output [7:0]  io_axi_ar_bits_len, // @[playground/src/cache/DCache.scala 83:14]
  output [2:0]  io_axi_ar_bits_size, // @[playground/src/cache/DCache.scala 83:14]
  output        io_axi_r_ready, // @[playground/src/cache/DCache.scala 83:14]
  input         io_axi_r_valid, // @[playground/src/cache/DCache.scala 83:14]
  input  [63:0] io_axi_r_bits_data, // @[playground/src/cache/DCache.scala 83:14]
  input  [1:0]  io_axi_r_bits_resp, // @[playground/src/cache/DCache.scala 83:14]
  input         io_axi_r_bits_last, // @[playground/src/cache/DCache.scala 83:14]
  input         io_axi_aw_ready, // @[playground/src/cache/DCache.scala 83:14]
  output        io_axi_aw_valid, // @[playground/src/cache/DCache.scala 83:14]
  output [31:0] io_axi_aw_bits_addr, // @[playground/src/cache/DCache.scala 83:14]
  output [7:0]  io_axi_aw_bits_len, // @[playground/src/cache/DCache.scala 83:14]
  output [2:0]  io_axi_aw_bits_size, // @[playground/src/cache/DCache.scala 83:14]
  input         io_axi_w_ready, // @[playground/src/cache/DCache.scala 83:14]
  output        io_axi_w_valid, // @[playground/src/cache/DCache.scala 83:14]
  output [63:0] io_axi_w_bits_data, // @[playground/src/cache/DCache.scala 83:14]
  output [7:0]  io_axi_w_bits_strb, // @[playground/src/cache/DCache.scala 83:14]
  output        io_axi_w_bits_last, // @[playground/src/cache/DCache.scala 83:14]
  output        io_axi_b_ready, // @[playground/src/cache/DCache.scala 83:14]
  input         io_axi_b_valid // @[playground/src/cache/DCache.scala 83:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [63:0] _RAND_333;
  reg [63:0] _RAND_334;
  reg [63:0] _RAND_335;
  reg [63:0] _RAND_336;
  reg [63:0] _RAND_337;
  reg [63:0] _RAND_338;
  reg [63:0] _RAND_339;
  reg [63:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [63:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [63:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
`endif // RANDOMIZE_REG_INIT
  wire  writeFifo_clock; // @[playground/src/cache/DCache.scala 151:34]
  wire  writeFifo_reset; // @[playground/src/cache/DCache.scala 151:34]
  wire  writeFifo_io_enq_ready; // @[playground/src/cache/DCache.scala 151:34]
  wire  writeFifo_io_enq_valid; // @[playground/src/cache/DCache.scala 151:34]
  wire [63:0] writeFifo_io_enq_bits_data; // @[playground/src/cache/DCache.scala 151:34]
  wire [63:0] writeFifo_io_enq_bits_addr; // @[playground/src/cache/DCache.scala 151:34]
  wire [7:0] writeFifo_io_enq_bits_strb; // @[playground/src/cache/DCache.scala 151:34]
  wire [2:0] writeFifo_io_enq_bits_size; // @[playground/src/cache/DCache.scala 151:34]
  wire  writeFifo_io_deq_ready; // @[playground/src/cache/DCache.scala 151:34]
  wire  writeFifo_io_deq_valid; // @[playground/src/cache/DCache.scala 151:34]
  wire [63:0] writeFifo_io_deq_bits_data; // @[playground/src/cache/DCache.scala 151:34]
  wire [63:0] writeFifo_io_deq_bits_addr; // @[playground/src/cache/DCache.scala 151:34]
  wire [7:0] writeFifo_io_deq_bits_strb; // @[playground/src/cache/DCache.scala 151:34]
  wire [2:0] writeFifo_io_deq_bits_size; // @[playground/src/cache/DCache.scala 151:34]
  wire  tagRam_0_clock; // @[playground/src/cache/DCache.scala 226:37]
  wire  tagRam_0_reset; // @[playground/src/cache/DCache.scala 226:37]
  wire [5:0] tagRam_0_io_raddr; // @[playground/src/cache/DCache.scala 226:37]
  wire [19:0] tagRam_0_io_rdata; // @[playground/src/cache/DCache.scala 226:37]
  wire [5:0] tagRam_0_io_waddr; // @[playground/src/cache/DCache.scala 226:37]
  wire [19:0] tagRam_0_io_wdata; // @[playground/src/cache/DCache.scala 226:37]
  wire  tagRam_0_io_wen; // @[playground/src/cache/DCache.scala 226:37]
  wire  tagRam_1_clock; // @[playground/src/cache/DCache.scala 226:37]
  wire  tagRam_1_reset; // @[playground/src/cache/DCache.scala 226:37]
  wire [5:0] tagRam_1_io_raddr; // @[playground/src/cache/DCache.scala 226:37]
  wire [19:0] tagRam_1_io_rdata; // @[playground/src/cache/DCache.scala 226:37]
  wire [5:0] tagRam_1_io_waddr; // @[playground/src/cache/DCache.scala 226:37]
  wire [19:0] tagRam_1_io_wdata; // @[playground/src/cache/DCache.scala 226:37]
  wire  tagRam_1_io_wen; // @[playground/src/cache/DCache.scala 226:37]
  wire  bank_0_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_0_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_0_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_0_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_0_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_0_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_0_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_0_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_2_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_2_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_2_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_2_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_2_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_2_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_2_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_2_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_3_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_3_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_3_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_3_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_3_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_3_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_3_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_3_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_4_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_4_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_4_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_4_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_4_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_4_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_4_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_4_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_5_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_5_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_5_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_5_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_5_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_5_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_5_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_5_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_6_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_6_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_6_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_6_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_6_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_6_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_6_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_6_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_7_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_7_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_7_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_7_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_7_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_7_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_7_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_7_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_0_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_0_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_0_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_0_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_0_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_0_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_0_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_0_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_1_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_1_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_1_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_1_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_1_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_1_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_1_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_1_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_2_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_2_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_2_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_2_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_2_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_2_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_2_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_2_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_3_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_3_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_3_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_3_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_3_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_3_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_3_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_3_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_4_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_4_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_4_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_4_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_4_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_4_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_4_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_4_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_5_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_5_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_5_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_5_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_5_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_5_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_5_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_5_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_6_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_6_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_6_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_6_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_6_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_6_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_6_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_6_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_7_1_clock; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_7_1_reset; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_7_1_io_raddr; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_7_1_io_rdata; // @[playground/src/cache/DCache.scala 228:38]
  wire [5:0] bank_7_1_io_waddr; // @[playground/src/cache/DCache.scala 228:38]
  wire  bank_7_1_io_wen; // @[playground/src/cache/DCache.scala 228:38]
  wire [7:0] bank_7_1_io_wstrb; // @[playground/src/cache/DCache.scala 228:38]
  wire [63:0] bank_7_1_io_wdata; // @[playground/src/cache/DCache.scala 228:38]
  reg [2:0] state; // @[playground/src/cache/DCache.scala 90:94]
  reg [2:0] ptw_state; // @[playground/src/cache/DCache.scala 94:103]
  wire  _ptw_working_T_1 = ptw_state != 3'h5; // @[playground/src/cache/DCache.scala 99:17]
  wire  _ptw_working_T_2 = ptw_state != 3'h0 & _ptw_working_T_1; // @[playground/src/cache/DCache.scala 98:33]
  wire  _ptw_working_T_4 = ~(io_cpu_tlb_ptw_pte_bits_access_fault | io_cpu_tlb_ptw_pte_bits_page_fault); // @[playground/src/cache/DCache.scala 100:7]
  wire  ptw_working = _ptw_working_T_2 & _ptw_working_T_4; // @[playground/src/cache/DCache.scala 99:29]
  reg [19:0] ptw_scratch_paddr_tag; // @[playground/src/cache/DCache.scala 101:28]
  reg [5:0] ptw_scratch_paddr_index; // @[playground/src/cache/DCache.scala 101:28]
  reg [5:0] ptw_scratch_paddr_offset; // @[playground/src/cache/DCache.scala 101:28]
  reg  ptw_scratch_replace; // @[playground/src/cache/DCache.scala 101:28]
  reg  ptw_scratch_dcache_wait; // @[playground/src/cache/DCache.scala 101:28]
  wire [5:0] exe_index = io_cpu_exe_addr[11:6]; // @[playground/src/cache/DCache.scala 117:34]
  wire [2:0] bank_index = io_cpu_addr[5:3]; // @[playground/src/cache/DCache.scala 119:31]
  reg  valid_0_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_0_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_1_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_1_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_2_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_2_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_3_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_3_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_4_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_4_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_5_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_5_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_6_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_6_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_7_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_7_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_8_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_8_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_9_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_9_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_10_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_10_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_11_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_11_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_12_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_12_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_13_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_13_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_14_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_14_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_15_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_15_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_16_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_16_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_17_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_17_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_18_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_18_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_19_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_19_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_20_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_20_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_21_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_21_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_22_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_22_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_23_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_23_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_24_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_24_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_25_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_25_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_26_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_26_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_27_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_27_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_28_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_28_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_29_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_29_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_30_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_30_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_31_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_31_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_32_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_32_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_33_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_33_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_34_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_34_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_35_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_35_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_36_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_36_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_37_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_37_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_38_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_38_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_39_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_39_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_40_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_40_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_41_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_41_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_42_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_42_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_43_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_43_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_44_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_44_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_45_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_45_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_46_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_46_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_47_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_47_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_48_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_48_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_49_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_49_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_50_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_50_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_51_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_51_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_52_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_52_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_53_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_53_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_54_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_54_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_55_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_55_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_56_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_56_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_57_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_57_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_58_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_58_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_59_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_59_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_60_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_60_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_61_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_61_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_62_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_62_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_63_0; // @[playground/src/cache/DCache.scala 134:22]
  reg  valid_63_1; // @[playground/src/cache/DCache.scala 134:22]
  reg  dirty_0_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_0_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_1_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_1_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_2_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_2_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_3_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_3_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_4_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_4_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_5_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_5_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_6_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_6_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_7_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_7_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_8_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_8_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_9_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_9_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_10_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_10_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_11_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_11_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_12_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_12_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_13_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_13_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_14_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_14_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_15_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_15_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_16_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_16_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_17_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_17_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_18_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_18_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_19_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_19_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_20_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_20_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_21_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_21_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_22_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_22_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_23_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_23_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_24_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_24_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_25_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_25_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_26_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_26_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_27_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_27_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_28_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_28_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_29_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_29_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_30_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_30_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_31_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_31_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_32_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_32_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_33_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_33_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_34_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_34_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_35_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_35_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_36_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_36_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_37_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_37_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_38_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_38_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_39_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_39_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_40_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_40_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_41_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_41_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_42_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_42_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_43_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_43_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_44_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_44_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_45_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_45_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_46_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_46_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_47_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_47_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_48_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_48_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_49_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_49_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_50_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_50_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_51_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_51_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_52_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_52_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_53_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_53_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_54_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_54_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_55_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_55_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_56_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_56_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_57_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_57_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_58_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_58_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_59_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_59_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_60_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_60_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_61_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_61_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_62_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_62_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_63_0; // @[playground/src/cache/DCache.scala 135:22]
  reg  dirty_63_1; // @[playground/src/cache/DCache.scala 135:22]
  reg  lru_0; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_1; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_2; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_3; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_4; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_5; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_6; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_7; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_8; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_9; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_10; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_11; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_12; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_13; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_14; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_15; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_16; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_17; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_18; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_19; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_20; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_21; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_22; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_23; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_24; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_25; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_26; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_27; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_28; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_29; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_30; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_31; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_32; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_33; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_34; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_35; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_36; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_37; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_38; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_39; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_40; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_41; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_42; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_43; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_44; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_45; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_46; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_47; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_48; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_49; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_50; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_51; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_52; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_53; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_54; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_55; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_56; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_57; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_58; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_59; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_60; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_61; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_62; // @[playground/src/cache/DCache.scala 136:22]
  reg  lru_63; // @[playground/src/cache/DCache.scala 136:22]
  wire [1:0] _dirty_index_T = {dirty_0_1,dirty_0_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_1 = |_dirty_index_T; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_2 = {dirty_1_1,dirty_1_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_3 = |_dirty_index_T_2; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_4 = {dirty_2_1,dirty_2_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_5 = |_dirty_index_T_4; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_6 = {dirty_3_1,dirty_3_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_7 = |_dirty_index_T_6; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_8 = {dirty_4_1,dirty_4_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_9 = |_dirty_index_T_8; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_10 = {dirty_5_1,dirty_5_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_11 = |_dirty_index_T_10; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_12 = {dirty_6_1,dirty_6_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_13 = |_dirty_index_T_12; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_14 = {dirty_7_1,dirty_7_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_15 = |_dirty_index_T_14; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_16 = {dirty_8_1,dirty_8_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_17 = |_dirty_index_T_16; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_18 = {dirty_9_1,dirty_9_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_19 = |_dirty_index_T_18; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_20 = {dirty_10_1,dirty_10_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_21 = |_dirty_index_T_20; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_22 = {dirty_11_1,dirty_11_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_23 = |_dirty_index_T_22; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_24 = {dirty_12_1,dirty_12_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_25 = |_dirty_index_T_24; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_26 = {dirty_13_1,dirty_13_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_27 = |_dirty_index_T_26; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_28 = {dirty_14_1,dirty_14_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_29 = |_dirty_index_T_28; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_30 = {dirty_15_1,dirty_15_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_31 = |_dirty_index_T_30; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_32 = {dirty_16_1,dirty_16_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_33 = |_dirty_index_T_32; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_34 = {dirty_17_1,dirty_17_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_35 = |_dirty_index_T_34; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_36 = {dirty_18_1,dirty_18_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_37 = |_dirty_index_T_36; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_38 = {dirty_19_1,dirty_19_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_39 = |_dirty_index_T_38; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_40 = {dirty_20_1,dirty_20_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_41 = |_dirty_index_T_40; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_42 = {dirty_21_1,dirty_21_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_43 = |_dirty_index_T_42; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_44 = {dirty_22_1,dirty_22_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_45 = |_dirty_index_T_44; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_46 = {dirty_23_1,dirty_23_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_47 = |_dirty_index_T_46; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_48 = {dirty_24_1,dirty_24_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_49 = |_dirty_index_T_48; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_50 = {dirty_25_1,dirty_25_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_51 = |_dirty_index_T_50; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_52 = {dirty_26_1,dirty_26_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_53 = |_dirty_index_T_52; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_54 = {dirty_27_1,dirty_27_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_55 = |_dirty_index_T_54; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_56 = {dirty_28_1,dirty_28_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_57 = |_dirty_index_T_56; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_58 = {dirty_29_1,dirty_29_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_59 = |_dirty_index_T_58; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_60 = {dirty_30_1,dirty_30_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_61 = |_dirty_index_T_60; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_62 = {dirty_31_1,dirty_31_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_63 = |_dirty_index_T_62; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_64 = {dirty_32_1,dirty_32_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_65 = |_dirty_index_T_64; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_66 = {dirty_33_1,dirty_33_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_67 = |_dirty_index_T_66; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_68 = {dirty_34_1,dirty_34_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_69 = |_dirty_index_T_68; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_70 = {dirty_35_1,dirty_35_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_71 = |_dirty_index_T_70; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_72 = {dirty_36_1,dirty_36_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_73 = |_dirty_index_T_72; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_74 = {dirty_37_1,dirty_37_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_75 = |_dirty_index_T_74; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_76 = {dirty_38_1,dirty_38_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_77 = |_dirty_index_T_76; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_78 = {dirty_39_1,dirty_39_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_79 = |_dirty_index_T_78; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_80 = {dirty_40_1,dirty_40_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_81 = |_dirty_index_T_80; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_82 = {dirty_41_1,dirty_41_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_83 = |_dirty_index_T_82; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_84 = {dirty_42_1,dirty_42_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_85 = |_dirty_index_T_84; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_86 = {dirty_43_1,dirty_43_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_87 = |_dirty_index_T_86; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_88 = {dirty_44_1,dirty_44_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_89 = |_dirty_index_T_88; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_90 = {dirty_45_1,dirty_45_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_91 = |_dirty_index_T_90; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_92 = {dirty_46_1,dirty_46_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_93 = |_dirty_index_T_92; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_94 = {dirty_47_1,dirty_47_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_95 = |_dirty_index_T_94; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_96 = {dirty_48_1,dirty_48_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_97 = |_dirty_index_T_96; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_98 = {dirty_49_1,dirty_49_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_99 = |_dirty_index_T_98; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_100 = {dirty_50_1,dirty_50_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_101 = |_dirty_index_T_100; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_102 = {dirty_51_1,dirty_51_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_103 = |_dirty_index_T_102; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_104 = {dirty_52_1,dirty_52_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_105 = |_dirty_index_T_104; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_106 = {dirty_53_1,dirty_53_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_107 = |_dirty_index_T_106; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_108 = {dirty_54_1,dirty_54_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_109 = |_dirty_index_T_108; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_110 = {dirty_55_1,dirty_55_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_111 = |_dirty_index_T_110; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_112 = {dirty_56_1,dirty_56_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_113 = |_dirty_index_T_112; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_114 = {dirty_57_1,dirty_57_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_115 = |_dirty_index_T_114; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_116 = {dirty_58_1,dirty_58_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_117 = |_dirty_index_T_116; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_118 = {dirty_59_1,dirty_59_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_119 = |_dirty_index_T_118; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_120 = {dirty_60_1,dirty_60_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_121 = |_dirty_index_T_120; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_122 = {dirty_61_1,dirty_61_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_123 = |_dirty_index_T_122; // @[playground/src/cache/DCache.scala 140:53]
  wire [1:0] _dirty_index_T_124 = {dirty_62_1,dirty_62_0}; // @[playground/src/cache/DCache.scala 140:46]
  wire  _dirty_index_T_125 = |_dirty_index_T_124; // @[playground/src/cache/DCache.scala 140:53]
  wire [5:0] _dirty_index_T_128 = _dirty_index_T_125 ? 6'h3e : 6'h3f; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_129 = _dirty_index_T_123 ? 6'h3d : _dirty_index_T_128; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_130 = _dirty_index_T_121 ? 6'h3c : _dirty_index_T_129; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_131 = _dirty_index_T_119 ? 6'h3b : _dirty_index_T_130; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_132 = _dirty_index_T_117 ? 6'h3a : _dirty_index_T_131; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_133 = _dirty_index_T_115 ? 6'h39 : _dirty_index_T_132; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_134 = _dirty_index_T_113 ? 6'h38 : _dirty_index_T_133; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_135 = _dirty_index_T_111 ? 6'h37 : _dirty_index_T_134; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_136 = _dirty_index_T_109 ? 6'h36 : _dirty_index_T_135; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_137 = _dirty_index_T_107 ? 6'h35 : _dirty_index_T_136; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_138 = _dirty_index_T_105 ? 6'h34 : _dirty_index_T_137; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_139 = _dirty_index_T_103 ? 6'h33 : _dirty_index_T_138; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_140 = _dirty_index_T_101 ? 6'h32 : _dirty_index_T_139; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_141 = _dirty_index_T_99 ? 6'h31 : _dirty_index_T_140; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_142 = _dirty_index_T_97 ? 6'h30 : _dirty_index_T_141; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_143 = _dirty_index_T_95 ? 6'h2f : _dirty_index_T_142; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_144 = _dirty_index_T_93 ? 6'h2e : _dirty_index_T_143; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_145 = _dirty_index_T_91 ? 6'h2d : _dirty_index_T_144; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_146 = _dirty_index_T_89 ? 6'h2c : _dirty_index_T_145; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_147 = _dirty_index_T_87 ? 6'h2b : _dirty_index_T_146; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_148 = _dirty_index_T_85 ? 6'h2a : _dirty_index_T_147; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_149 = _dirty_index_T_83 ? 6'h29 : _dirty_index_T_148; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_150 = _dirty_index_T_81 ? 6'h28 : _dirty_index_T_149; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_151 = _dirty_index_T_79 ? 6'h27 : _dirty_index_T_150; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_152 = _dirty_index_T_77 ? 6'h26 : _dirty_index_T_151; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_153 = _dirty_index_T_75 ? 6'h25 : _dirty_index_T_152; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_154 = _dirty_index_T_73 ? 6'h24 : _dirty_index_T_153; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_155 = _dirty_index_T_71 ? 6'h23 : _dirty_index_T_154; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_156 = _dirty_index_T_69 ? 6'h22 : _dirty_index_T_155; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_157 = _dirty_index_T_67 ? 6'h21 : _dirty_index_T_156; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_158 = _dirty_index_T_65 ? 6'h20 : _dirty_index_T_157; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_159 = _dirty_index_T_63 ? 6'h1f : _dirty_index_T_158; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_160 = _dirty_index_T_61 ? 6'h1e : _dirty_index_T_159; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_161 = _dirty_index_T_59 ? 6'h1d : _dirty_index_T_160; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_162 = _dirty_index_T_57 ? 6'h1c : _dirty_index_T_161; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_163 = _dirty_index_T_55 ? 6'h1b : _dirty_index_T_162; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_164 = _dirty_index_T_53 ? 6'h1a : _dirty_index_T_163; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_165 = _dirty_index_T_51 ? 6'h19 : _dirty_index_T_164; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_166 = _dirty_index_T_49 ? 6'h18 : _dirty_index_T_165; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_167 = _dirty_index_T_47 ? 6'h17 : _dirty_index_T_166; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_168 = _dirty_index_T_45 ? 6'h16 : _dirty_index_T_167; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_169 = _dirty_index_T_43 ? 6'h15 : _dirty_index_T_168; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_170 = _dirty_index_T_41 ? 6'h14 : _dirty_index_T_169; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_171 = _dirty_index_T_39 ? 6'h13 : _dirty_index_T_170; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_172 = _dirty_index_T_37 ? 6'h12 : _dirty_index_T_171; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_173 = _dirty_index_T_35 ? 6'h11 : _dirty_index_T_172; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_174 = _dirty_index_T_33 ? 6'h10 : _dirty_index_T_173; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_175 = _dirty_index_T_31 ? 6'hf : _dirty_index_T_174; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_176 = _dirty_index_T_29 ? 6'he : _dirty_index_T_175; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_177 = _dirty_index_T_27 ? 6'hd : _dirty_index_T_176; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_178 = _dirty_index_T_25 ? 6'hc : _dirty_index_T_177; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_179 = _dirty_index_T_23 ? 6'hb : _dirty_index_T_178; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_180 = _dirty_index_T_21 ? 6'ha : _dirty_index_T_179; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_181 = _dirty_index_T_19 ? 6'h9 : _dirty_index_T_180; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_182 = _dirty_index_T_17 ? 6'h8 : _dirty_index_T_181; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_183 = _dirty_index_T_15 ? 6'h7 : _dirty_index_T_182; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_184 = _dirty_index_T_13 ? 6'h6 : _dirty_index_T_183; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_185 = _dirty_index_T_11 ? 6'h5 : _dirty_index_T_184; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_186 = _dirty_index_T_9 ? 6'h4 : _dirty_index_T_185; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_187 = _dirty_index_T_7 ? 6'h3 : _dirty_index_T_186; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_188 = _dirty_index_T_5 ? 6'h2 : _dirty_index_T_187; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _dirty_index_T_189 = _dirty_index_T_3 ? 6'h1 : _dirty_index_T_188; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] dirty_index = _dirty_index_T_1 ? 6'h0 : _dirty_index_T_189; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  reg  fence; // @[playground/src/cache/DCache.scala 145:22]
  reg  readsram; // @[playground/src/cache/DCache.scala 148:25]
  reg  writeFifo_axi_busy; // @[playground/src/cache/DCache.scala 152:35]
  reg [7:0] burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22]
  reg [7:0] burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22]
  reg [2:0] bank_wbindex; // @[playground/src/cache/DCache.scala 165:29]
  reg [63:0] bank_wbdata_0; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_1; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_2; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_3; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_4; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_5; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_6; // @[playground/src/cache/DCache.scala 166:29]
  reg [63:0] bank_wbdata_7; // @[playground/src/cache/DCache.scala 166:29]
  wire  _use_next_addr_T = state == 3'h0; // @[playground/src/cache/DCache.scala 169:30]
  wire  _use_next_addr_T_1 = state == 3'h4; // @[playground/src/cache/DCache.scala 169:52]
  wire  use_next_addr = state == 3'h0 | state == 3'h4; // @[playground/src/cache/DCache.scala 169:42]
  reg  do_replace; // @[playground/src/cache/DCache.scala 170:30]
  reg [19:0] ppn; // @[playground/src/cache/DCache.scala 567:28]
  reg [1:0] vpn_index; // @[playground/src/cache/DCache.scala 568:28]
  wire  _vpnn_T = vpn_index == 2'h0; // @[playground/src/cache/DCache.scala 615:22]
  wire [8:0] vpn_vpn0 = io_cpu_tlb_ptw_vpn_bits[8:0]; // @[playground/src/cache/DCache.scala 565:53]
  wire [8:0] _vpnn_T_3 = _vpnn_T ? vpn_vpn0 : 9'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _vpnn_T_1 = vpn_index == 2'h1; // @[playground/src/cache/DCache.scala 616:22]
  wire [8:0] vpn_vpn1 = io_cpu_tlb_ptw_vpn_bits[17:9]; // @[playground/src/cache/DCache.scala 565:53]
  wire [8:0] _vpnn_T_4 = _vpnn_T_1 ? vpn_vpn1 : 9'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [8:0] _vpnn_T_6 = _vpnn_T_3 | _vpnn_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _vpnn_T_2 = vpn_index == 2'h2; // @[playground/src/cache/DCache.scala 617:22]
  wire [8:0] vpn_vpn2 = io_cpu_tlb_ptw_vpn_bits[26:18]; // @[playground/src/cache/DCache.scala 565:53]
  wire [8:0] _vpnn_T_5 = _vpnn_T_2 ? vpn_vpn2 : 9'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [8:0] vpnn = _vpnn_T_6 | _vpnn_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _ptw_addr_T_1 = {ppn,vpnn,3'h0}; // @[playground/src/defines/TlbBundles.scala 58:8]
  wire [19:0] ptw_addr_tag = _ptw_addr_T_1[31:12]; // @[playground/src/cache/DCache.scala 620:56]
  wire [5:0] ptw_addr_index = _ptw_addr_T_1[11:6]; // @[playground/src/cache/DCache.scala 620:56]
  wire [5:0] ptw_addr_offset = _ptw_addr_T_1[5:0]; // @[playground/src/cache/DCache.scala 620:56]
  wire [31:0] _pte_uncached_T = {ptw_addr_tag,ptw_addr_index,ptw_addr_offset}; // @[playground/src/cache/DCache.scala 621:55]
  wire [31:0] _pte_uncached_T_1 = _pte_uncached_T ^ 32'h30000000; // @[playground/src/defines/Const.scala 78:13]
  wire  _pte_uncached_T_3 = _pte_uncached_T_1[31:28] == 4'h0; // @[playground/src/defines/Const.scala 78:48]
  wire [31:0] _pte_uncached_T_4 = _pte_uncached_T ^ 32'h40000000; // @[playground/src/defines/Const.scala 78:13]
  wire  _pte_uncached_T_6 = _pte_uncached_T_4[31:30] == 2'h0; // @[playground/src/defines/Const.scala 78:48]
  wire  pte_uncached = _pte_uncached_T_3 | _pte_uncached_T_6; // @[playground/src/defines/Const.scala 80:15]
  wire [5:0] _GEN_5427 = pte_uncached ? io_cpu_addr[11:6] : ptw_addr_index; // @[playground/src/cache/DCache.scala 173:17 622:26 632:31]
  wire [5:0] _GEN_5841 = 3'h2 == ptw_state ? ptw_scratch_paddr_index : io_cpu_addr[11:6]; // @[playground/src/cache/DCache.scala 173:17 603:21 641:29]
  wire [5:0] _GEN_5884 = 3'h1 == ptw_state ? _GEN_5427 : _GEN_5841; // @[playground/src/cache/DCache.scala 603:21]
  wire [5:0] replace_index = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  wire [5:0] tag_rindex = use_next_addr ? exe_index : replace_index; // @[playground/src/cache/DCache.scala 181:23]
  reg  tag_wstrb_0; // @[playground/src/cache/DCache.scala 182:27]
  reg  tag_wstrb_1; // @[playground/src/cache/DCache.scala 182:27]
  reg [19:0] tag_wdata; // @[playground/src/cache/DCache.scala 183:27]
  reg [19:0] tag_0; // @[playground/src/cache/DCache.scala 187:20]
  reg [19:0] tag_1; // @[playground/src/cache/DCache.scala 187:20]
  wire  _GEN_145 = 6'h1 == replace_index ? valid_1_0 : valid_0_0; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_146 = 6'h2 == replace_index ? valid_2_0 : _GEN_145; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_147 = 6'h3 == replace_index ? valid_3_0 : _GEN_146; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_148 = 6'h4 == replace_index ? valid_4_0 : _GEN_147; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_149 = 6'h5 == replace_index ? valid_5_0 : _GEN_148; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_150 = 6'h6 == replace_index ? valid_6_0 : _GEN_149; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_151 = 6'h7 == replace_index ? valid_7_0 : _GEN_150; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_152 = 6'h8 == replace_index ? valid_8_0 : _GEN_151; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_153 = 6'h9 == replace_index ? valid_9_0 : _GEN_152; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_154 = 6'ha == replace_index ? valid_10_0 : _GEN_153; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_155 = 6'hb == replace_index ? valid_11_0 : _GEN_154; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_156 = 6'hc == replace_index ? valid_12_0 : _GEN_155; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_157 = 6'hd == replace_index ? valid_13_0 : _GEN_156; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_158 = 6'he == replace_index ? valid_14_0 : _GEN_157; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_159 = 6'hf == replace_index ? valid_15_0 : _GEN_158; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_160 = 6'h10 == replace_index ? valid_16_0 : _GEN_159; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_161 = 6'h11 == replace_index ? valid_17_0 : _GEN_160; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_162 = 6'h12 == replace_index ? valid_18_0 : _GEN_161; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_163 = 6'h13 == replace_index ? valid_19_0 : _GEN_162; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_164 = 6'h14 == replace_index ? valid_20_0 : _GEN_163; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_165 = 6'h15 == replace_index ? valid_21_0 : _GEN_164; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_166 = 6'h16 == replace_index ? valid_22_0 : _GEN_165; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_167 = 6'h17 == replace_index ? valid_23_0 : _GEN_166; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_168 = 6'h18 == replace_index ? valid_24_0 : _GEN_167; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_169 = 6'h19 == replace_index ? valid_25_0 : _GEN_168; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_170 = 6'h1a == replace_index ? valid_26_0 : _GEN_169; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_171 = 6'h1b == replace_index ? valid_27_0 : _GEN_170; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_172 = 6'h1c == replace_index ? valid_28_0 : _GEN_171; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_173 = 6'h1d == replace_index ? valid_29_0 : _GEN_172; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_174 = 6'h1e == replace_index ? valid_30_0 : _GEN_173; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_175 = 6'h1f == replace_index ? valid_31_0 : _GEN_174; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_176 = 6'h20 == replace_index ? valid_32_0 : _GEN_175; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_177 = 6'h21 == replace_index ? valid_33_0 : _GEN_176; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_178 = 6'h22 == replace_index ? valid_34_0 : _GEN_177; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_179 = 6'h23 == replace_index ? valid_35_0 : _GEN_178; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_180 = 6'h24 == replace_index ? valid_36_0 : _GEN_179; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_181 = 6'h25 == replace_index ? valid_37_0 : _GEN_180; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_182 = 6'h26 == replace_index ? valid_38_0 : _GEN_181; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_183 = 6'h27 == replace_index ? valid_39_0 : _GEN_182; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_184 = 6'h28 == replace_index ? valid_40_0 : _GEN_183; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_185 = 6'h29 == replace_index ? valid_41_0 : _GEN_184; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_186 = 6'h2a == replace_index ? valid_42_0 : _GEN_185; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_187 = 6'h2b == replace_index ? valid_43_0 : _GEN_186; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_188 = 6'h2c == replace_index ? valid_44_0 : _GEN_187; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_189 = 6'h2d == replace_index ? valid_45_0 : _GEN_188; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_190 = 6'h2e == replace_index ? valid_46_0 : _GEN_189; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_191 = 6'h2f == replace_index ? valid_47_0 : _GEN_190; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_192 = 6'h30 == replace_index ? valid_48_0 : _GEN_191; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_193 = 6'h31 == replace_index ? valid_49_0 : _GEN_192; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_194 = 6'h32 == replace_index ? valid_50_0 : _GEN_193; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_195 = 6'h33 == replace_index ? valid_51_0 : _GEN_194; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_196 = 6'h34 == replace_index ? valid_52_0 : _GEN_195; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_197 = 6'h35 == replace_index ? valid_53_0 : _GEN_196; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_198 = 6'h36 == replace_index ? valid_54_0 : _GEN_197; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_199 = 6'h37 == replace_index ? valid_55_0 : _GEN_198; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_200 = 6'h38 == replace_index ? valid_56_0 : _GEN_199; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_201 = 6'h39 == replace_index ? valid_57_0 : _GEN_200; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_202 = 6'h3a == replace_index ? valid_58_0 : _GEN_201; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_203 = 6'h3b == replace_index ? valid_59_0 : _GEN_202; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_204 = 6'h3c == replace_index ? valid_60_0 : _GEN_203; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_205 = 6'h3d == replace_index ? valid_61_0 : _GEN_204; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_206 = 6'h3e == replace_index ? valid_62_0 : _GEN_205; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_207 = 6'h3f == replace_index ? valid_63_0 : _GEN_206; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _tag_compare_valid_0_T_22 = tag_0 == io_cpu_tlb_ptag & _GEN_207; // @[playground/src/cache/DCache.scala 247:36]
  wire  _tag_compare_valid_0_T_23 = _tag_compare_valid_0_T_22 & io_cpu_tlb_hit; // @[playground/src/cache/DCache.scala 248:33]
  wire  _GEN_5433 = 6'h1 == ptw_scratch_paddr_index ? valid_1_0 : valid_0_0; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5434 = 6'h2 == ptw_scratch_paddr_index ? valid_2_0 : _GEN_5433; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5435 = 6'h3 == ptw_scratch_paddr_index ? valid_3_0 : _GEN_5434; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5436 = 6'h4 == ptw_scratch_paddr_index ? valid_4_0 : _GEN_5435; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5437 = 6'h5 == ptw_scratch_paddr_index ? valid_5_0 : _GEN_5436; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5438 = 6'h6 == ptw_scratch_paddr_index ? valid_6_0 : _GEN_5437; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5439 = 6'h7 == ptw_scratch_paddr_index ? valid_7_0 : _GEN_5438; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5440 = 6'h8 == ptw_scratch_paddr_index ? valid_8_0 : _GEN_5439; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5441 = 6'h9 == ptw_scratch_paddr_index ? valid_9_0 : _GEN_5440; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5442 = 6'ha == ptw_scratch_paddr_index ? valid_10_0 : _GEN_5441; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5443 = 6'hb == ptw_scratch_paddr_index ? valid_11_0 : _GEN_5442; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5444 = 6'hc == ptw_scratch_paddr_index ? valid_12_0 : _GEN_5443; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5445 = 6'hd == ptw_scratch_paddr_index ? valid_13_0 : _GEN_5444; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5446 = 6'he == ptw_scratch_paddr_index ? valid_14_0 : _GEN_5445; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5447 = 6'hf == ptw_scratch_paddr_index ? valid_15_0 : _GEN_5446; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5448 = 6'h10 == ptw_scratch_paddr_index ? valid_16_0 : _GEN_5447; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5449 = 6'h11 == ptw_scratch_paddr_index ? valid_17_0 : _GEN_5448; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5450 = 6'h12 == ptw_scratch_paddr_index ? valid_18_0 : _GEN_5449; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5451 = 6'h13 == ptw_scratch_paddr_index ? valid_19_0 : _GEN_5450; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5452 = 6'h14 == ptw_scratch_paddr_index ? valid_20_0 : _GEN_5451; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5453 = 6'h15 == ptw_scratch_paddr_index ? valid_21_0 : _GEN_5452; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5454 = 6'h16 == ptw_scratch_paddr_index ? valid_22_0 : _GEN_5453; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5455 = 6'h17 == ptw_scratch_paddr_index ? valid_23_0 : _GEN_5454; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5456 = 6'h18 == ptw_scratch_paddr_index ? valid_24_0 : _GEN_5455; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5457 = 6'h19 == ptw_scratch_paddr_index ? valid_25_0 : _GEN_5456; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5458 = 6'h1a == ptw_scratch_paddr_index ? valid_26_0 : _GEN_5457; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5459 = 6'h1b == ptw_scratch_paddr_index ? valid_27_0 : _GEN_5458; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5460 = 6'h1c == ptw_scratch_paddr_index ? valid_28_0 : _GEN_5459; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5461 = 6'h1d == ptw_scratch_paddr_index ? valid_29_0 : _GEN_5460; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5462 = 6'h1e == ptw_scratch_paddr_index ? valid_30_0 : _GEN_5461; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5463 = 6'h1f == ptw_scratch_paddr_index ? valid_31_0 : _GEN_5462; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5464 = 6'h20 == ptw_scratch_paddr_index ? valid_32_0 : _GEN_5463; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5465 = 6'h21 == ptw_scratch_paddr_index ? valid_33_0 : _GEN_5464; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5466 = 6'h22 == ptw_scratch_paddr_index ? valid_34_0 : _GEN_5465; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5467 = 6'h23 == ptw_scratch_paddr_index ? valid_35_0 : _GEN_5466; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5468 = 6'h24 == ptw_scratch_paddr_index ? valid_36_0 : _GEN_5467; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5469 = 6'h25 == ptw_scratch_paddr_index ? valid_37_0 : _GEN_5468; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5470 = 6'h26 == ptw_scratch_paddr_index ? valid_38_0 : _GEN_5469; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5471 = 6'h27 == ptw_scratch_paddr_index ? valid_39_0 : _GEN_5470; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5472 = 6'h28 == ptw_scratch_paddr_index ? valid_40_0 : _GEN_5471; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5473 = 6'h29 == ptw_scratch_paddr_index ? valid_41_0 : _GEN_5472; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5474 = 6'h2a == ptw_scratch_paddr_index ? valid_42_0 : _GEN_5473; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5475 = 6'h2b == ptw_scratch_paddr_index ? valid_43_0 : _GEN_5474; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5476 = 6'h2c == ptw_scratch_paddr_index ? valid_44_0 : _GEN_5475; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5477 = 6'h2d == ptw_scratch_paddr_index ? valid_45_0 : _GEN_5476; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5478 = 6'h2e == ptw_scratch_paddr_index ? valid_46_0 : _GEN_5477; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5479 = 6'h2f == ptw_scratch_paddr_index ? valid_47_0 : _GEN_5478; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5480 = 6'h30 == ptw_scratch_paddr_index ? valid_48_0 : _GEN_5479; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5481 = 6'h31 == ptw_scratch_paddr_index ? valid_49_0 : _GEN_5480; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5482 = 6'h32 == ptw_scratch_paddr_index ? valid_50_0 : _GEN_5481; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5483 = 6'h33 == ptw_scratch_paddr_index ? valid_51_0 : _GEN_5482; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5484 = 6'h34 == ptw_scratch_paddr_index ? valid_52_0 : _GEN_5483; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5485 = 6'h35 == ptw_scratch_paddr_index ? valid_53_0 : _GEN_5484; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5486 = 6'h36 == ptw_scratch_paddr_index ? valid_54_0 : _GEN_5485; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5487 = 6'h37 == ptw_scratch_paddr_index ? valid_55_0 : _GEN_5486; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5488 = 6'h38 == ptw_scratch_paddr_index ? valid_56_0 : _GEN_5487; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5489 = 6'h39 == ptw_scratch_paddr_index ? valid_57_0 : _GEN_5488; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5490 = 6'h3a == ptw_scratch_paddr_index ? valid_58_0 : _GEN_5489; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5491 = 6'h3b == ptw_scratch_paddr_index ? valid_59_0 : _GEN_5490; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5492 = 6'h3c == ptw_scratch_paddr_index ? valid_60_0 : _GEN_5491; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5493 = 6'h3d == ptw_scratch_paddr_index ? valid_61_0 : _GEN_5492; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5494 = 6'h3e == ptw_scratch_paddr_index ? valid_62_0 : _GEN_5493; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5495 = 6'h3f == ptw_scratch_paddr_index ? valid_63_0 : _GEN_5494; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _tag_compare_valid_0_T_25 = tag_0 == ptw_scratch_paddr_tag & _GEN_5495; // @[playground/src/cache/DCache.scala 644:44]
  wire  _GEN_5842 = 3'h2 == ptw_state ? _tag_compare_valid_0_T_25 : _tag_compare_valid_0_T_23; // @[playground/src/cache/DCache.scala 603:21 246:28 643:30]
  wire  _GEN_5889 = 3'h1 == ptw_state ? _tag_compare_valid_0_T_23 : _GEN_5842; // @[playground/src/cache/DCache.scala 603:21 246:28]
  wire  tag_compare_valid_0 = 3'h0 == ptw_state ? _tag_compare_valid_0_T_23 : _GEN_5889; // @[playground/src/cache/DCache.scala 603:21 246:28]
  wire  _GEN_209 = 6'h1 == replace_index ? valid_1_1 : valid_0_1; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_210 = 6'h2 == replace_index ? valid_2_1 : _GEN_209; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_211 = 6'h3 == replace_index ? valid_3_1 : _GEN_210; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_212 = 6'h4 == replace_index ? valid_4_1 : _GEN_211; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_213 = 6'h5 == replace_index ? valid_5_1 : _GEN_212; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_214 = 6'h6 == replace_index ? valid_6_1 : _GEN_213; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_215 = 6'h7 == replace_index ? valid_7_1 : _GEN_214; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_216 = 6'h8 == replace_index ? valid_8_1 : _GEN_215; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_217 = 6'h9 == replace_index ? valid_9_1 : _GEN_216; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_218 = 6'ha == replace_index ? valid_10_1 : _GEN_217; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_219 = 6'hb == replace_index ? valid_11_1 : _GEN_218; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_220 = 6'hc == replace_index ? valid_12_1 : _GEN_219; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_221 = 6'hd == replace_index ? valid_13_1 : _GEN_220; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_222 = 6'he == replace_index ? valid_14_1 : _GEN_221; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_223 = 6'hf == replace_index ? valid_15_1 : _GEN_222; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_224 = 6'h10 == replace_index ? valid_16_1 : _GEN_223; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_225 = 6'h11 == replace_index ? valid_17_1 : _GEN_224; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_226 = 6'h12 == replace_index ? valid_18_1 : _GEN_225; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_227 = 6'h13 == replace_index ? valid_19_1 : _GEN_226; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_228 = 6'h14 == replace_index ? valid_20_1 : _GEN_227; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_229 = 6'h15 == replace_index ? valid_21_1 : _GEN_228; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_230 = 6'h16 == replace_index ? valid_22_1 : _GEN_229; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_231 = 6'h17 == replace_index ? valid_23_1 : _GEN_230; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_232 = 6'h18 == replace_index ? valid_24_1 : _GEN_231; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_233 = 6'h19 == replace_index ? valid_25_1 : _GEN_232; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_234 = 6'h1a == replace_index ? valid_26_1 : _GEN_233; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_235 = 6'h1b == replace_index ? valid_27_1 : _GEN_234; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_236 = 6'h1c == replace_index ? valid_28_1 : _GEN_235; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_237 = 6'h1d == replace_index ? valid_29_1 : _GEN_236; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_238 = 6'h1e == replace_index ? valid_30_1 : _GEN_237; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_239 = 6'h1f == replace_index ? valid_31_1 : _GEN_238; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_240 = 6'h20 == replace_index ? valid_32_1 : _GEN_239; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_241 = 6'h21 == replace_index ? valid_33_1 : _GEN_240; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_242 = 6'h22 == replace_index ? valid_34_1 : _GEN_241; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_243 = 6'h23 == replace_index ? valid_35_1 : _GEN_242; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_244 = 6'h24 == replace_index ? valid_36_1 : _GEN_243; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_245 = 6'h25 == replace_index ? valid_37_1 : _GEN_244; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_246 = 6'h26 == replace_index ? valid_38_1 : _GEN_245; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_247 = 6'h27 == replace_index ? valid_39_1 : _GEN_246; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_248 = 6'h28 == replace_index ? valid_40_1 : _GEN_247; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_249 = 6'h29 == replace_index ? valid_41_1 : _GEN_248; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_250 = 6'h2a == replace_index ? valid_42_1 : _GEN_249; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_251 = 6'h2b == replace_index ? valid_43_1 : _GEN_250; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_252 = 6'h2c == replace_index ? valid_44_1 : _GEN_251; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_253 = 6'h2d == replace_index ? valid_45_1 : _GEN_252; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_254 = 6'h2e == replace_index ? valid_46_1 : _GEN_253; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_255 = 6'h2f == replace_index ? valid_47_1 : _GEN_254; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_256 = 6'h30 == replace_index ? valid_48_1 : _GEN_255; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_257 = 6'h31 == replace_index ? valid_49_1 : _GEN_256; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_258 = 6'h32 == replace_index ? valid_50_1 : _GEN_257; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_259 = 6'h33 == replace_index ? valid_51_1 : _GEN_258; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_260 = 6'h34 == replace_index ? valid_52_1 : _GEN_259; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_261 = 6'h35 == replace_index ? valid_53_1 : _GEN_260; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_262 = 6'h36 == replace_index ? valid_54_1 : _GEN_261; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_263 = 6'h37 == replace_index ? valid_55_1 : _GEN_262; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_264 = 6'h38 == replace_index ? valid_56_1 : _GEN_263; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_265 = 6'h39 == replace_index ? valid_57_1 : _GEN_264; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_266 = 6'h3a == replace_index ? valid_58_1 : _GEN_265; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_267 = 6'h3b == replace_index ? valid_59_1 : _GEN_266; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_268 = 6'h3c == replace_index ? valid_60_1 : _GEN_267; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_269 = 6'h3d == replace_index ? valid_61_1 : _GEN_268; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_270 = 6'h3e == replace_index ? valid_62_1 : _GEN_269; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _GEN_271 = 6'h3f == replace_index ? valid_63_1 : _GEN_270; // @[playground/src/cache/DCache.scala 247:{36,36}]
  wire  _tag_compare_valid_1_T_22 = tag_1 == io_cpu_tlb_ptag & _GEN_271; // @[playground/src/cache/DCache.scala 247:36]
  wire  _tag_compare_valid_1_T_23 = _tag_compare_valid_1_T_22 & io_cpu_tlb_hit; // @[playground/src/cache/DCache.scala 248:33]
  wire  _GEN_5497 = 6'h1 == ptw_scratch_paddr_index ? valid_1_1 : valid_0_1; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5498 = 6'h2 == ptw_scratch_paddr_index ? valid_2_1 : _GEN_5497; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5499 = 6'h3 == ptw_scratch_paddr_index ? valid_3_1 : _GEN_5498; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5500 = 6'h4 == ptw_scratch_paddr_index ? valid_4_1 : _GEN_5499; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5501 = 6'h5 == ptw_scratch_paddr_index ? valid_5_1 : _GEN_5500; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5502 = 6'h6 == ptw_scratch_paddr_index ? valid_6_1 : _GEN_5501; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5503 = 6'h7 == ptw_scratch_paddr_index ? valid_7_1 : _GEN_5502; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5504 = 6'h8 == ptw_scratch_paddr_index ? valid_8_1 : _GEN_5503; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5505 = 6'h9 == ptw_scratch_paddr_index ? valid_9_1 : _GEN_5504; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5506 = 6'ha == ptw_scratch_paddr_index ? valid_10_1 : _GEN_5505; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5507 = 6'hb == ptw_scratch_paddr_index ? valid_11_1 : _GEN_5506; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5508 = 6'hc == ptw_scratch_paddr_index ? valid_12_1 : _GEN_5507; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5509 = 6'hd == ptw_scratch_paddr_index ? valid_13_1 : _GEN_5508; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5510 = 6'he == ptw_scratch_paddr_index ? valid_14_1 : _GEN_5509; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5511 = 6'hf == ptw_scratch_paddr_index ? valid_15_1 : _GEN_5510; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5512 = 6'h10 == ptw_scratch_paddr_index ? valid_16_1 : _GEN_5511; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5513 = 6'h11 == ptw_scratch_paddr_index ? valid_17_1 : _GEN_5512; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5514 = 6'h12 == ptw_scratch_paddr_index ? valid_18_1 : _GEN_5513; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5515 = 6'h13 == ptw_scratch_paddr_index ? valid_19_1 : _GEN_5514; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5516 = 6'h14 == ptw_scratch_paddr_index ? valid_20_1 : _GEN_5515; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5517 = 6'h15 == ptw_scratch_paddr_index ? valid_21_1 : _GEN_5516; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5518 = 6'h16 == ptw_scratch_paddr_index ? valid_22_1 : _GEN_5517; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5519 = 6'h17 == ptw_scratch_paddr_index ? valid_23_1 : _GEN_5518; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5520 = 6'h18 == ptw_scratch_paddr_index ? valid_24_1 : _GEN_5519; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5521 = 6'h19 == ptw_scratch_paddr_index ? valid_25_1 : _GEN_5520; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5522 = 6'h1a == ptw_scratch_paddr_index ? valid_26_1 : _GEN_5521; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5523 = 6'h1b == ptw_scratch_paddr_index ? valid_27_1 : _GEN_5522; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5524 = 6'h1c == ptw_scratch_paddr_index ? valid_28_1 : _GEN_5523; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5525 = 6'h1d == ptw_scratch_paddr_index ? valid_29_1 : _GEN_5524; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5526 = 6'h1e == ptw_scratch_paddr_index ? valid_30_1 : _GEN_5525; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5527 = 6'h1f == ptw_scratch_paddr_index ? valid_31_1 : _GEN_5526; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5528 = 6'h20 == ptw_scratch_paddr_index ? valid_32_1 : _GEN_5527; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5529 = 6'h21 == ptw_scratch_paddr_index ? valid_33_1 : _GEN_5528; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5530 = 6'h22 == ptw_scratch_paddr_index ? valid_34_1 : _GEN_5529; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5531 = 6'h23 == ptw_scratch_paddr_index ? valid_35_1 : _GEN_5530; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5532 = 6'h24 == ptw_scratch_paddr_index ? valid_36_1 : _GEN_5531; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5533 = 6'h25 == ptw_scratch_paddr_index ? valid_37_1 : _GEN_5532; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5534 = 6'h26 == ptw_scratch_paddr_index ? valid_38_1 : _GEN_5533; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5535 = 6'h27 == ptw_scratch_paddr_index ? valid_39_1 : _GEN_5534; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5536 = 6'h28 == ptw_scratch_paddr_index ? valid_40_1 : _GEN_5535; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5537 = 6'h29 == ptw_scratch_paddr_index ? valid_41_1 : _GEN_5536; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5538 = 6'h2a == ptw_scratch_paddr_index ? valid_42_1 : _GEN_5537; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5539 = 6'h2b == ptw_scratch_paddr_index ? valid_43_1 : _GEN_5538; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5540 = 6'h2c == ptw_scratch_paddr_index ? valid_44_1 : _GEN_5539; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5541 = 6'h2d == ptw_scratch_paddr_index ? valid_45_1 : _GEN_5540; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5542 = 6'h2e == ptw_scratch_paddr_index ? valid_46_1 : _GEN_5541; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5543 = 6'h2f == ptw_scratch_paddr_index ? valid_47_1 : _GEN_5542; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5544 = 6'h30 == ptw_scratch_paddr_index ? valid_48_1 : _GEN_5543; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5545 = 6'h31 == ptw_scratch_paddr_index ? valid_49_1 : _GEN_5544; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5546 = 6'h32 == ptw_scratch_paddr_index ? valid_50_1 : _GEN_5545; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5547 = 6'h33 == ptw_scratch_paddr_index ? valid_51_1 : _GEN_5546; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5548 = 6'h34 == ptw_scratch_paddr_index ? valid_52_1 : _GEN_5547; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5549 = 6'h35 == ptw_scratch_paddr_index ? valid_53_1 : _GEN_5548; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5550 = 6'h36 == ptw_scratch_paddr_index ? valid_54_1 : _GEN_5549; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5551 = 6'h37 == ptw_scratch_paddr_index ? valid_55_1 : _GEN_5550; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5552 = 6'h38 == ptw_scratch_paddr_index ? valid_56_1 : _GEN_5551; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5553 = 6'h39 == ptw_scratch_paddr_index ? valid_57_1 : _GEN_5552; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5554 = 6'h3a == ptw_scratch_paddr_index ? valid_58_1 : _GEN_5553; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5555 = 6'h3b == ptw_scratch_paddr_index ? valid_59_1 : _GEN_5554; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5556 = 6'h3c == ptw_scratch_paddr_index ? valid_60_1 : _GEN_5555; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5557 = 6'h3d == ptw_scratch_paddr_index ? valid_61_1 : _GEN_5556; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5558 = 6'h3e == ptw_scratch_paddr_index ? valid_62_1 : _GEN_5557; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _GEN_5559 = 6'h3f == ptw_scratch_paddr_index ? valid_63_1 : _GEN_5558; // @[playground/src/cache/DCache.scala 644:{44,44}]
  wire  _tag_compare_valid_1_T_25 = tag_1 == ptw_scratch_paddr_tag & _GEN_5559; // @[playground/src/cache/DCache.scala 644:44]
  wire  _GEN_5843 = 3'h2 == ptw_state ? _tag_compare_valid_1_T_25 : _tag_compare_valid_1_T_23; // @[playground/src/cache/DCache.scala 603:21 246:28 643:30]
  wire  _GEN_5890 = 3'h1 == ptw_state ? _tag_compare_valid_1_T_23 : _GEN_5843; // @[playground/src/cache/DCache.scala 603:21 246:28]
  wire  tag_compare_valid_1 = 3'h0 == ptw_state ? _tag_compare_valid_1_T_23 : _GEN_5890; // @[playground/src/cache/DCache.scala 603:21 246:28]
  wire  cache_hit = tag_compare_valid_0 | tag_compare_valid_1; // @[playground/src/cache/DCache.scala 190:53]
  wire  _mmio_read_stall_T = |io_cpu_wen; // @[playground/src/cache/DCache.scala 192:61]
  wire  mmio_read_stall = io_cpu_tlb_uncached & ~(|io_cpu_wen); // @[playground/src/cache/DCache.scala 192:46]
  wire  mmio_write_stall = io_cpu_tlb_uncached & _mmio_read_stall_T & ~writeFifo_io_enq_ready; // @[playground/src/cache/DCache.scala 193:64]
  wire  _cached_stall_T = ~io_cpu_tlb_uncached; // @[playground/src/cache/DCache.scala 194:26]
  wire  _cached_stall_T_1 = ~cache_hit; // @[playground/src/cache/DCache.scala 194:50]
  wire  cached_stall = ~io_cpu_tlb_uncached & ~cache_hit; // @[playground/src/cache/DCache.scala 194:47]
  wire  _dcache_stall_T_3 = ~io_cpu_tlb_hit; // @[playground/src/cache/DCache.scala 202:63]
  wire  _dcache_stall_T_4 = cached_stall | mmio_read_stall | mmio_write_stall | ~io_cpu_tlb_hit; // @[playground/src/cache/DCache.scala 202:60]
  wire  _dcache_stall_T_5 = io_cpu_fence_i | fence; // @[playground/src/cache/DCache.scala 203:22]
  wire  _dcache_stall_T_6 = io_cpu_en ? _dcache_stall_T_4 : _dcache_stall_T_5; // @[playground/src/cache/DCache.scala 200:8]
  wire  _dcache_stall_T_7 = state != 3'h4; // @[playground/src/cache/DCache.scala 205:11]
  wire  dcache_stall = _use_next_addr_T ? _dcache_stall_T_6 : _dcache_stall_T_7; // @[playground/src/cache/DCache.scala 198:25]
  wire  _io_cpu_dcache_ready_T = ~dcache_stall; // @[playground/src/cache/DCache.scala 207:26]
  reg [63:0] saved_rdata; // @[playground/src/cache/DCache.scala 209:28]
  wire [63:0] data_0_0 = bank_0_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] data_0_1 = bank_0_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5962 = 3'h0 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_1 = 3'h0 == bank_index & tag_compare_valid_1 ? data_0_1 : data_0_0; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_1_0 = bank_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5963 = 3'h1 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire  _GEN_5964 = ~tag_compare_valid_1; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_2 = 3'h1 == bank_index & ~tag_compare_valid_1 ? data_1_0 : _GEN_1; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_1_1 = bank_1_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_3 = 3'h1 == bank_index & tag_compare_valid_1 ? data_1_1 : _GEN_2; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_2_0 = bank_2_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5966 = 3'h2 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_4 = 3'h2 == bank_index & ~tag_compare_valid_1 ? data_2_0 : _GEN_3; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_2_1 = bank_2_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_5 = 3'h2 == bank_index & tag_compare_valid_1 ? data_2_1 : _GEN_4; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_3_0 = bank_3_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5969 = 3'h3 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_6 = 3'h3 == bank_index & ~tag_compare_valid_1 ? data_3_0 : _GEN_5; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_3_1 = bank_3_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_7 = 3'h3 == bank_index & tag_compare_valid_1 ? data_3_1 : _GEN_6; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_4_0 = bank_4_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5972 = 3'h4 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_8 = 3'h4 == bank_index & ~tag_compare_valid_1 ? data_4_0 : _GEN_7; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_4_1 = bank_4_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_9 = 3'h4 == bank_index & tag_compare_valid_1 ? data_4_1 : _GEN_8; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_5_0 = bank_5_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5975 = 3'h5 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_10 = 3'h5 == bank_index & ~tag_compare_valid_1 ? data_5_0 : _GEN_9; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_5_1 = bank_5_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_11 = 3'h5 == bank_index & tag_compare_valid_1 ? data_5_1 : _GEN_10; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_6_0 = bank_6_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5978 = 3'h6 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_12 = 3'h6 == bank_index & ~tag_compare_valid_1 ? data_6_0 : _GEN_11; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_6_1 = bank_6_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_13 = 3'h6 == bank_index & tag_compare_valid_1 ? data_6_1 : _GEN_12; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_7_0 = bank_7_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire  _GEN_5981 = 3'h7 == bank_index; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] _GEN_14 = 3'h7 == bank_index & ~tag_compare_valid_1 ? data_7_0 : _GEN_13; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [63:0] data_7_1 = bank_7_1_io_rdata; // @[playground/src/cache/DCache.scala 185:18 232:24]
  wire [63:0] _GEN_15 = 3'h7 == bank_index & tag_compare_valid_1 ? data_7_1 : _GEN_14; // @[playground/src/cache/DCache.scala 211:{22,22}]
  wire [5:0] _bank_raddr_T_2 = state == 3'h2 ? dirty_index : tag_rindex; // @[playground/src/cache/DCache.scala 218:20]
  wire [7:0] wstrb_0_0 = _GEN_5962 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_0_1 = _GEN_5962 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_1_0 = _GEN_5963 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_1_1 = _GEN_5963 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_2_0 = _GEN_5966 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_2_1 = _GEN_5966 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_3_0 = _GEN_5969 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_3_1 = _GEN_5969 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_4_0 = _GEN_5972 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_4_1 = _GEN_5972 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_5_0 = _GEN_5975 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_5_1 = _GEN_5975 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_6_0 = _GEN_5978 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_6_1 = _GEN_5978 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_7_0 = _GEN_5981 & _GEN_5964 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire [7:0] wstrb_7_1 = _GEN_5981 & tag_compare_valid_1 ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 222:33 223:{33,33}]
  wire  _replace_wstrb_0_0_T_6 = tag_compare_valid_0 & io_cpu_en & _mmio_read_stall_T & _cached_stall_T &
    _use_next_addr_T; // @[playground/src/cache/DCache.scala 252:85]
  wire [7:0] _replace_wstrb_0_0_T_9 = burst_wstrb_0[0] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_0_0 = _replace_wstrb_0_0_T_6 ? wstrb_0_0 : _replace_wstrb_0_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_1_0_T_9 = burst_wstrb_0[1] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_1_0 = _replace_wstrb_0_0_T_6 ? wstrb_1_0 : _replace_wstrb_1_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_2_0_T_9 = burst_wstrb_0[2] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_2_0 = _replace_wstrb_0_0_T_6 ? wstrb_2_0 : _replace_wstrb_2_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_3_0_T_9 = burst_wstrb_0[3] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_3_0 = _replace_wstrb_0_0_T_6 ? wstrb_3_0 : _replace_wstrb_3_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_4_0_T_9 = burst_wstrb_0[4] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_4_0 = _replace_wstrb_0_0_T_6 ? wstrb_4_0 : _replace_wstrb_4_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_5_0_T_9 = burst_wstrb_0[5] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_5_0 = _replace_wstrb_0_0_T_6 ? wstrb_5_0 : _replace_wstrb_5_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_6_0_T_9 = burst_wstrb_0[6] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_6_0 = _replace_wstrb_0_0_T_6 ? wstrb_6_0 : _replace_wstrb_6_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_7_0_T_9 = burst_wstrb_0[7] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_7_0 = _replace_wstrb_0_0_T_6 ? wstrb_7_0 : _replace_wstrb_7_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire  _replace_wstrb_0_1_T_6 = tag_compare_valid_1 & io_cpu_en & _mmio_read_stall_T & _cached_stall_T &
    _use_next_addr_T; // @[playground/src/cache/DCache.scala 252:85]
  wire [7:0] _replace_wstrb_0_1_T_9 = burst_wstrb_1[0] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_0_1 = _replace_wstrb_0_1_T_6 ? wstrb_0_1 : _replace_wstrb_0_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_1_1_T_9 = burst_wstrb_1[1] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_1_1 = _replace_wstrb_0_1_T_6 ? wstrb_1_1 : _replace_wstrb_1_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_2_1_T_9 = burst_wstrb_1[2] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_2_1 = _replace_wstrb_0_1_T_6 ? wstrb_2_1 : _replace_wstrb_2_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_3_1_T_9 = burst_wstrb_1[3] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_3_1 = _replace_wstrb_0_1_T_6 ? wstrb_3_1 : _replace_wstrb_3_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_4_1_T_9 = burst_wstrb_1[4] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_4_1 = _replace_wstrb_0_1_T_6 ? wstrb_4_1 : _replace_wstrb_4_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_5_1_T_9 = burst_wstrb_1[5] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_5_1 = _replace_wstrb_0_1_T_6 ? wstrb_5_1 : _replace_wstrb_5_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_6_1_T_9 = burst_wstrb_1[6] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_6_1 = _replace_wstrb_0_1_T_6 ? wstrb_6_1 : _replace_wstrb_6_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  wire [7:0] _replace_wstrb_7_1_T_9 = burst_wstrb_1[7] ? 8'hff : 8'h0; // @[playground/src/cache/DCache.scala 254:13]
  wire [7:0] replace_wstrb_7_1 = _replace_wstrb_0_1_T_6 ? wstrb_7_1 : _replace_wstrb_7_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  reg [31:0] ar_addr; // @[playground/src/cache/DCache.scala 259:24]
  reg [7:0] ar_len; // @[playground/src/cache/DCache.scala 259:24]
  reg [2:0] ar_size; // @[playground/src/cache/DCache.scala 259:24]
  reg  arvalid; // @[playground/src/cache/DCache.scala 260:24]
  reg  rready; // @[playground/src/cache/DCache.scala 263:23]
  reg [31:0] aw_addr; // @[playground/src/cache/DCache.scala 265:24]
  reg [7:0] aw_len; // @[playground/src/cache/DCache.scala 265:24]
  reg [2:0] aw_size; // @[playground/src/cache/DCache.scala 265:24]
  reg  awvalid; // @[playground/src/cache/DCache.scala 266:24]
  reg [63:0] w_data; // @[playground/src/cache/DCache.scala 269:23]
  reg [7:0] w_strb; // @[playground/src/cache/DCache.scala 269:23]
  reg  w_last; // @[playground/src/cache/DCache.scala 269:23]
  reg  wvalid; // @[playground/src/cache/DCache.scala 270:23]
  reg  access_fault; // @[playground/src/cache/DCache.scala 277:29]
  reg  page_fault; // @[playground/src/cache/DCache.scala 278:29]
  wire  _addr_err_T_27 = io_cpu_addr[39] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_29 = io_cpu_addr[40] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_31 = io_cpu_addr[41] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_33 = io_cpu_addr[42] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_35 = io_cpu_addr[43] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_37 = io_cpu_addr[44] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_39 = io_cpu_addr[45] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_41 = io_cpu_addr[46] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_43 = io_cpu_addr[47] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_45 = io_cpu_addr[48] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_47 = io_cpu_addr[49] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_49 = io_cpu_addr[50] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_51 = io_cpu_addr[51] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_53 = io_cpu_addr[52] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_55 = io_cpu_addr[53] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_57 = io_cpu_addr[54] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_59 = io_cpu_addr[55] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_61 = io_cpu_addr[56] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_63 = io_cpu_addr[57] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_65 = io_cpu_addr[58] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_67 = io_cpu_addr[59] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_69 = io_cpu_addr[60] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_71 = io_cpu_addr[61] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_73 = io_cpu_addr[62] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  _addr_err_T_75 = io_cpu_addr[63] != io_cpu_addr[38]; // @[playground/src/cache/DCache.scala 283:12]
  wire  addr_err = _addr_err_T_27 | _addr_err_T_29 | _addr_err_T_31 | _addr_err_T_33 | _addr_err_T_35 | _addr_err_T_37
     | _addr_err_T_39 | _addr_err_T_41 | _addr_err_T_43 | _addr_err_T_45 | _addr_err_T_47 | _addr_err_T_49 |
    _addr_err_T_51 | _addr_err_T_53 | _addr_err_T_55 | _addr_err_T_57 | _addr_err_T_59 | _addr_err_T_61 | _addr_err_T_63
     | _addr_err_T_65 | _addr_err_T_67 | _addr_err_T_69 | _addr_err_T_71 | _addr_err_T_73 | _addr_err_T_75; // @[playground/src/cache/DCache.scala 284:15]
  wire  _T = io_axi_aw_ready & io_axi_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _GEN_272 = _T ? 1'h0 : awvalid; // @[playground/src/cache/DCache.scala 291:26 292:15 266:24]
  wire  _T_1 = io_axi_w_ready & io_axi_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _GEN_273 = _T_1 ? 1'h0 : wvalid; // @[playground/src/cache/DCache.scala 294:25 295:14 270:23]
  wire  _GEN_274 = _T_1 ? 1'h0 : w_last; // @[playground/src/cache/DCache.scala 294:25 296:14 269:23]
  wire  _T_2 = io_axi_b_ready & io_axi_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_3 = writeFifo_io_deq_ready & writeFifo_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [63:0] _GEN_276 = _T_3 ? writeFifo_io_deq_bits_addr : {{32'd0}, aw_addr}; // @[playground/src/cache/DCache.scala 303:33 304:15 265:24]
  wire [2:0] _GEN_277 = _T_3 ? writeFifo_io_deq_bits_size : aw_size; // @[playground/src/cache/DCache.scala 303:33 305:15 265:24]
  wire [63:0] _GEN_278 = _T_3 ? writeFifo_io_deq_bits_data : w_data; // @[playground/src/cache/DCache.scala 303:33 306:15 269:23]
  wire [7:0] _GEN_279 = _T_3 ? writeFifo_io_deq_bits_strb : w_strb; // @[playground/src/cache/DCache.scala 303:33 307:15 269:23]
  wire  _GEN_280 = writeFifo_io_deq_valid; // @[playground/src/cache/DCache.scala 157:26 301:38 302:28]
  wire [63:0] _GEN_281 = writeFifo_io_deq_valid ? _GEN_276 : {{32'd0}, aw_addr}; // @[playground/src/cache/DCache.scala 265:24 301:38]
  wire [2:0] _GEN_282 = writeFifo_io_deq_valid ? _GEN_277 : aw_size; // @[playground/src/cache/DCache.scala 265:24 301:38]
  wire [63:0] _GEN_283 = writeFifo_io_deq_valid ? _GEN_278 : w_data; // @[playground/src/cache/DCache.scala 269:23 301:38]
  wire [7:0] _GEN_284 = writeFifo_io_deq_valid ? _GEN_279 : w_strb; // @[playground/src/cache/DCache.scala 269:23 301:38]
  wire [7:0] _GEN_285 = writeFifo_io_deq_valid ? 8'h0 : aw_len; // @[playground/src/cache/DCache.scala 265:24 301:38 309:24]
  wire  _GEN_286 = writeFifo_io_deq_valid | awvalid; // @[playground/src/cache/DCache.scala 266:24 301:38 310:24]
  wire  _GEN_287 = writeFifo_io_deq_valid | w_last; // @[playground/src/cache/DCache.scala 269:23 301:38 311:24]
  wire  _GEN_288 = writeFifo_io_deq_valid | wvalid; // @[playground/src/cache/DCache.scala 270:23 301:38 312:24]
  wire  _GEN_289 = writeFifo_io_deq_valid | writeFifo_axi_busy; // @[playground/src/cache/DCache.scala 301:38 313:24 152:35]
  wire  _GEN_290 = writeFifo_axi_busy ? _GEN_272 : _GEN_286; // @[playground/src/cache/DCache.scala 290:28]
  wire  _GEN_291 = writeFifo_axi_busy ? _GEN_273 : _GEN_288; // @[playground/src/cache/DCache.scala 290:28]
  wire  _GEN_292 = writeFifo_axi_busy ? _GEN_274 : _GEN_287; // @[playground/src/cache/DCache.scala 290:28]
  wire [63:0] _GEN_295 = writeFifo_axi_busy ? {{32'd0}, aw_addr} : _GEN_281; // @[playground/src/cache/DCache.scala 265:24 290:28]
  wire [2:0] _GEN_296 = writeFifo_axi_busy ? aw_size : _GEN_282; // @[playground/src/cache/DCache.scala 265:24 290:28]
  wire [63:0] _GEN_297 = writeFifo_axi_busy ? w_data : _GEN_283; // @[playground/src/cache/DCache.scala 269:23 290:28]
  wire [7:0] _GEN_298 = writeFifo_axi_busy ? w_strb : _GEN_284; // @[playground/src/cache/DCache.scala 269:23 290:28]
  wire [7:0] _GEN_299 = writeFifo_axi_busy ? aw_len : _GEN_285; // @[playground/src/cache/DCache.scala 265:24 290:28]
  wire  _T_7 = ~io_cpu_complete_single_request; // @[playground/src/cache/DCache.scala 334:20]
  wire [2:0] _GEN_300 = ~io_cpu_complete_single_request ? 3'h4 : state; // @[playground/src/cache/DCache.scala 334:53 335:23 90:94]
  wire  _GEN_301 = writeFifo_io_enq_ready; // @[playground/src/cache/DCache.scala 155:26 327:42 328:42]
  wire [63:0] _GEN_302 = writeFifo_io_enq_ready ? {{32'd0}, io_cpu_tlb_paddr} : 64'h0; // @[playground/src/cache/DCache.scala 156:26 327:42 329:42]
  wire [7:0] _GEN_303 = writeFifo_io_enq_ready ? io_cpu_rlen : 8'h0; // @[playground/src/cache/DCache.scala 156:26 327:42 330:42]
  wire [7:0] _GEN_304 = writeFifo_io_enq_ready ? io_cpu_wstrb : 8'h0; // @[playground/src/cache/DCache.scala 156:26 327:42 331:42]
  wire [63:0] _GEN_305 = writeFifo_io_enq_ready ? io_cpu_wdata : 64'h0; // @[playground/src/cache/DCache.scala 156:26 327:42 332:42]
  wire [2:0] _GEN_306 = writeFifo_io_enq_ready ? _GEN_300 : state; // @[playground/src/cache/DCache.scala 327:42 90:94]
  wire  _T_8 = ~writeFifo_io_deq_valid; // @[playground/src/cache/DCache.scala 338:22]
  wire [31:0] _GEN_307 = ~writeFifo_io_deq_valid ? io_cpu_tlb_paddr : ar_addr; // @[playground/src/cache/DCache.scala 338:39 339:21 259:24]
  wire [7:0] _GEN_308 = ~writeFifo_io_deq_valid ? 8'h0 : ar_len; // @[playground/src/cache/DCache.scala 338:39 340:21 259:24]
  wire [7:0] _GEN_309 = ~writeFifo_io_deq_valid ? io_cpu_rlen : {{5'd0}, ar_size}; // @[playground/src/cache/DCache.scala 338:39 341:21 259:24]
  wire  _GEN_310 = ~writeFifo_io_deq_valid | arvalid; // @[playground/src/cache/DCache.scala 338:39 342:21 260:24]
  wire [2:0] _GEN_311 = ~writeFifo_io_deq_valid ? 3'h1 : state; // @[playground/src/cache/DCache.scala 338:39 343:21 90:94]
  wire  _GEN_312 = ~writeFifo_io_deq_valid | rready; // @[playground/src/cache/DCache.scala 338:39 344:21 263:23]
  wire  _GEN_313 = _mmio_read_stall_T & _GEN_301; // @[playground/src/cache/DCache.scala 155:26 326:32]
  wire [63:0] _GEN_314 = _mmio_read_stall_T ? _GEN_302 : 64'h0; // @[playground/src/cache/DCache.scala 156:26 326:32]
  wire [7:0] _GEN_315 = _mmio_read_stall_T ? _GEN_303 : 8'h0; // @[playground/src/cache/DCache.scala 156:26 326:32]
  wire [7:0] _GEN_316 = _mmio_read_stall_T ? _GEN_304 : 8'h0; // @[playground/src/cache/DCache.scala 156:26 326:32]
  wire [63:0] _GEN_317 = _mmio_read_stall_T ? _GEN_305 : 64'h0; // @[playground/src/cache/DCache.scala 156:26 326:32]
  wire [2:0] _GEN_318 = _mmio_read_stall_T ? _GEN_306 : _GEN_311; // @[playground/src/cache/DCache.scala 326:32]
  wire [31:0] _GEN_319 = _mmio_read_stall_T ? ar_addr : _GEN_307; // @[playground/src/cache/DCache.scala 259:24 326:32]
  wire [7:0] _GEN_320 = _mmio_read_stall_T ? ar_len : _GEN_308; // @[playground/src/cache/DCache.scala 259:24 326:32]
  wire [7:0] _GEN_321 = _mmio_read_stall_T ? {{5'd0}, ar_size} : _GEN_309; // @[playground/src/cache/DCache.scala 259:24 326:32]
  wire  _GEN_322 = _mmio_read_stall_T ? arvalid : _GEN_310; // @[playground/src/cache/DCache.scala 260:24 326:32]
  wire  _GEN_323 = _mmio_read_stall_T ? rready : _GEN_312; // @[playground/src/cache/DCache.scala 263:23 326:32]
  wire  _GEN_324 = 6'h0 == replace_index ? _GEN_5964 : lru_0; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_325 = 6'h1 == replace_index ? _GEN_5964 : lru_1; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_326 = 6'h2 == replace_index ? _GEN_5964 : lru_2; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_327 = 6'h3 == replace_index ? _GEN_5964 : lru_3; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_328 = 6'h4 == replace_index ? _GEN_5964 : lru_4; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_329 = 6'h5 == replace_index ? _GEN_5964 : lru_5; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_330 = 6'h6 == replace_index ? _GEN_5964 : lru_6; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_331 = 6'h7 == replace_index ? _GEN_5964 : lru_7; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_332 = 6'h8 == replace_index ? _GEN_5964 : lru_8; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_333 = 6'h9 == replace_index ? _GEN_5964 : lru_9; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_334 = 6'ha == replace_index ? _GEN_5964 : lru_10; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_335 = 6'hb == replace_index ? _GEN_5964 : lru_11; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_336 = 6'hc == replace_index ? _GEN_5964 : lru_12; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_337 = 6'hd == replace_index ? _GEN_5964 : lru_13; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_338 = 6'he == replace_index ? _GEN_5964 : lru_14; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_339 = 6'hf == replace_index ? _GEN_5964 : lru_15; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_340 = 6'h10 == replace_index ? _GEN_5964 : lru_16; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_341 = 6'h11 == replace_index ? _GEN_5964 : lru_17; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_342 = 6'h12 == replace_index ? _GEN_5964 : lru_18; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_343 = 6'h13 == replace_index ? _GEN_5964 : lru_19; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_344 = 6'h14 == replace_index ? _GEN_5964 : lru_20; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_345 = 6'h15 == replace_index ? _GEN_5964 : lru_21; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_346 = 6'h16 == replace_index ? _GEN_5964 : lru_22; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_347 = 6'h17 == replace_index ? _GEN_5964 : lru_23; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_348 = 6'h18 == replace_index ? _GEN_5964 : lru_24; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_349 = 6'h19 == replace_index ? _GEN_5964 : lru_25; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_350 = 6'h1a == replace_index ? _GEN_5964 : lru_26; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_351 = 6'h1b == replace_index ? _GEN_5964 : lru_27; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_352 = 6'h1c == replace_index ? _GEN_5964 : lru_28; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_353 = 6'h1d == replace_index ? _GEN_5964 : lru_29; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_354 = 6'h1e == replace_index ? _GEN_5964 : lru_30; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_355 = 6'h1f == replace_index ? _GEN_5964 : lru_31; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_356 = 6'h20 == replace_index ? _GEN_5964 : lru_32; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_357 = 6'h21 == replace_index ? _GEN_5964 : lru_33; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_358 = 6'h22 == replace_index ? _GEN_5964 : lru_34; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_359 = 6'h23 == replace_index ? _GEN_5964 : lru_35; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_360 = 6'h24 == replace_index ? _GEN_5964 : lru_36; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_361 = 6'h25 == replace_index ? _GEN_5964 : lru_37; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_362 = 6'h26 == replace_index ? _GEN_5964 : lru_38; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_363 = 6'h27 == replace_index ? _GEN_5964 : lru_39; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_364 = 6'h28 == replace_index ? _GEN_5964 : lru_40; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_365 = 6'h29 == replace_index ? _GEN_5964 : lru_41; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_366 = 6'h2a == replace_index ? _GEN_5964 : lru_42; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_367 = 6'h2b == replace_index ? _GEN_5964 : lru_43; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_368 = 6'h2c == replace_index ? _GEN_5964 : lru_44; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_369 = 6'h2d == replace_index ? _GEN_5964 : lru_45; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_370 = 6'h2e == replace_index ? _GEN_5964 : lru_46; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_371 = 6'h2f == replace_index ? _GEN_5964 : lru_47; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_372 = 6'h30 == replace_index ? _GEN_5964 : lru_48; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_373 = 6'h31 == replace_index ? _GEN_5964 : lru_49; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_374 = 6'h32 == replace_index ? _GEN_5964 : lru_50; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_375 = 6'h33 == replace_index ? _GEN_5964 : lru_51; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_376 = 6'h34 == replace_index ? _GEN_5964 : lru_52; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_377 = 6'h35 == replace_index ? _GEN_5964 : lru_53; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_378 = 6'h36 == replace_index ? _GEN_5964 : lru_54; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_379 = 6'h37 == replace_index ? _GEN_5964 : lru_55; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_380 = 6'h38 == replace_index ? _GEN_5964 : lru_56; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_381 = 6'h39 == replace_index ? _GEN_5964 : lru_57; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_382 = 6'h3a == replace_index ? _GEN_5964 : lru_58; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_383 = 6'h3b == replace_index ? _GEN_5964 : lru_59; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_384 = 6'h3c == replace_index ? _GEN_5964 : lru_60; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_385 = 6'h3d == replace_index ? _GEN_5964 : lru_61; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_386 = 6'h3e == replace_index ? _GEN_5964 : lru_62; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_387 = 6'h3f == replace_index ? _GEN_5964 : lru_63; // @[playground/src/cache/DCache.scala 136:22 352:{27,27}]
  wire  _GEN_6288 = 6'h0 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_388 = 6'h0 == replace_index & _GEN_5964 | dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_389 = 6'h0 == replace_index & tag_compare_valid_1 | dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6293 = 6'h1 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_390 = 6'h1 == replace_index & _GEN_5964 | dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_391 = 6'h1 == replace_index & tag_compare_valid_1 | dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6298 = 6'h2 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_392 = 6'h2 == replace_index & _GEN_5964 | dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_393 = 6'h2 == replace_index & tag_compare_valid_1 | dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6303 = 6'h3 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_394 = 6'h3 == replace_index & _GEN_5964 | dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_395 = 6'h3 == replace_index & tag_compare_valid_1 | dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6308 = 6'h4 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_396 = 6'h4 == replace_index & _GEN_5964 | dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_397 = 6'h4 == replace_index & tag_compare_valid_1 | dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6313 = 6'h5 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_398 = 6'h5 == replace_index & _GEN_5964 | dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_399 = 6'h5 == replace_index & tag_compare_valid_1 | dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6318 = 6'h6 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_400 = 6'h6 == replace_index & _GEN_5964 | dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_401 = 6'h6 == replace_index & tag_compare_valid_1 | dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6323 = 6'h7 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_402 = 6'h7 == replace_index & _GEN_5964 | dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_403 = 6'h7 == replace_index & tag_compare_valid_1 | dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6328 = 6'h8 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_404 = 6'h8 == replace_index & _GEN_5964 | dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_405 = 6'h8 == replace_index & tag_compare_valid_1 | dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6333 = 6'h9 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_406 = 6'h9 == replace_index & _GEN_5964 | dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_407 = 6'h9 == replace_index & tag_compare_valid_1 | dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6338 = 6'ha == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_408 = 6'ha == replace_index & _GEN_5964 | dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_409 = 6'ha == replace_index & tag_compare_valid_1 | dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6343 = 6'hb == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_410 = 6'hb == replace_index & _GEN_5964 | dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_411 = 6'hb == replace_index & tag_compare_valid_1 | dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6348 = 6'hc == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_412 = 6'hc == replace_index & _GEN_5964 | dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_413 = 6'hc == replace_index & tag_compare_valid_1 | dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6353 = 6'hd == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_414 = 6'hd == replace_index & _GEN_5964 | dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_415 = 6'hd == replace_index & tag_compare_valid_1 | dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6358 = 6'he == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_416 = 6'he == replace_index & _GEN_5964 | dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_417 = 6'he == replace_index & tag_compare_valid_1 | dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6363 = 6'hf == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_418 = 6'hf == replace_index & _GEN_5964 | dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_419 = 6'hf == replace_index & tag_compare_valid_1 | dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6368 = 6'h10 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_420 = 6'h10 == replace_index & _GEN_5964 | dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_421 = 6'h10 == replace_index & tag_compare_valid_1 | dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6373 = 6'h11 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_422 = 6'h11 == replace_index & _GEN_5964 | dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_423 = 6'h11 == replace_index & tag_compare_valid_1 | dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6378 = 6'h12 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_424 = 6'h12 == replace_index & _GEN_5964 | dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_425 = 6'h12 == replace_index & tag_compare_valid_1 | dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6383 = 6'h13 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_426 = 6'h13 == replace_index & _GEN_5964 | dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_427 = 6'h13 == replace_index & tag_compare_valid_1 | dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6388 = 6'h14 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_428 = 6'h14 == replace_index & _GEN_5964 | dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_429 = 6'h14 == replace_index & tag_compare_valid_1 | dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6393 = 6'h15 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_430 = 6'h15 == replace_index & _GEN_5964 | dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_431 = 6'h15 == replace_index & tag_compare_valid_1 | dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6398 = 6'h16 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_432 = 6'h16 == replace_index & _GEN_5964 | dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_433 = 6'h16 == replace_index & tag_compare_valid_1 | dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6403 = 6'h17 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_434 = 6'h17 == replace_index & _GEN_5964 | dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_435 = 6'h17 == replace_index & tag_compare_valid_1 | dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6408 = 6'h18 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_436 = 6'h18 == replace_index & _GEN_5964 | dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_437 = 6'h18 == replace_index & tag_compare_valid_1 | dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6413 = 6'h19 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_438 = 6'h19 == replace_index & _GEN_5964 | dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_439 = 6'h19 == replace_index & tag_compare_valid_1 | dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6418 = 6'h1a == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_440 = 6'h1a == replace_index & _GEN_5964 | dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_441 = 6'h1a == replace_index & tag_compare_valid_1 | dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6423 = 6'h1b == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_442 = 6'h1b == replace_index & _GEN_5964 | dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_443 = 6'h1b == replace_index & tag_compare_valid_1 | dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6428 = 6'h1c == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_444 = 6'h1c == replace_index & _GEN_5964 | dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_445 = 6'h1c == replace_index & tag_compare_valid_1 | dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6433 = 6'h1d == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_446 = 6'h1d == replace_index & _GEN_5964 | dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_447 = 6'h1d == replace_index & tag_compare_valid_1 | dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6438 = 6'h1e == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_448 = 6'h1e == replace_index & _GEN_5964 | dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_449 = 6'h1e == replace_index & tag_compare_valid_1 | dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6443 = 6'h1f == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_450 = 6'h1f == replace_index & _GEN_5964 | dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_451 = 6'h1f == replace_index & tag_compare_valid_1 | dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6448 = 6'h20 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_452 = 6'h20 == replace_index & _GEN_5964 | dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_453 = 6'h20 == replace_index & tag_compare_valid_1 | dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6453 = 6'h21 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_454 = 6'h21 == replace_index & _GEN_5964 | dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_455 = 6'h21 == replace_index & tag_compare_valid_1 | dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6458 = 6'h22 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_456 = 6'h22 == replace_index & _GEN_5964 | dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_457 = 6'h22 == replace_index & tag_compare_valid_1 | dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6463 = 6'h23 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_458 = 6'h23 == replace_index & _GEN_5964 | dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_459 = 6'h23 == replace_index & tag_compare_valid_1 | dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6468 = 6'h24 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_460 = 6'h24 == replace_index & _GEN_5964 | dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_461 = 6'h24 == replace_index & tag_compare_valid_1 | dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6473 = 6'h25 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_462 = 6'h25 == replace_index & _GEN_5964 | dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_463 = 6'h25 == replace_index & tag_compare_valid_1 | dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6478 = 6'h26 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_464 = 6'h26 == replace_index & _GEN_5964 | dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_465 = 6'h26 == replace_index & tag_compare_valid_1 | dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6483 = 6'h27 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_466 = 6'h27 == replace_index & _GEN_5964 | dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_467 = 6'h27 == replace_index & tag_compare_valid_1 | dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6488 = 6'h28 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_468 = 6'h28 == replace_index & _GEN_5964 | dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_469 = 6'h28 == replace_index & tag_compare_valid_1 | dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6493 = 6'h29 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_470 = 6'h29 == replace_index & _GEN_5964 | dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_471 = 6'h29 == replace_index & tag_compare_valid_1 | dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6498 = 6'h2a == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_472 = 6'h2a == replace_index & _GEN_5964 | dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_473 = 6'h2a == replace_index & tag_compare_valid_1 | dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6503 = 6'h2b == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_474 = 6'h2b == replace_index & _GEN_5964 | dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_475 = 6'h2b == replace_index & tag_compare_valid_1 | dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6508 = 6'h2c == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_476 = 6'h2c == replace_index & _GEN_5964 | dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_477 = 6'h2c == replace_index & tag_compare_valid_1 | dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6513 = 6'h2d == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_478 = 6'h2d == replace_index & _GEN_5964 | dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_479 = 6'h2d == replace_index & tag_compare_valid_1 | dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6518 = 6'h2e == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_480 = 6'h2e == replace_index & _GEN_5964 | dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_481 = 6'h2e == replace_index & tag_compare_valid_1 | dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6523 = 6'h2f == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_482 = 6'h2f == replace_index & _GEN_5964 | dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_483 = 6'h2f == replace_index & tag_compare_valid_1 | dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6528 = 6'h30 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_484 = 6'h30 == replace_index & _GEN_5964 | dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_485 = 6'h30 == replace_index & tag_compare_valid_1 | dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6533 = 6'h31 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_486 = 6'h31 == replace_index & _GEN_5964 | dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_487 = 6'h31 == replace_index & tag_compare_valid_1 | dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6538 = 6'h32 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_488 = 6'h32 == replace_index & _GEN_5964 | dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_489 = 6'h32 == replace_index & tag_compare_valid_1 | dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6543 = 6'h33 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_490 = 6'h33 == replace_index & _GEN_5964 | dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_491 = 6'h33 == replace_index & tag_compare_valid_1 | dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6548 = 6'h34 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_492 = 6'h34 == replace_index & _GEN_5964 | dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_493 = 6'h34 == replace_index & tag_compare_valid_1 | dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6553 = 6'h35 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_494 = 6'h35 == replace_index & _GEN_5964 | dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_495 = 6'h35 == replace_index & tag_compare_valid_1 | dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6558 = 6'h36 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_496 = 6'h36 == replace_index & _GEN_5964 | dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_497 = 6'h36 == replace_index & tag_compare_valid_1 | dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6563 = 6'h37 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_498 = 6'h37 == replace_index & _GEN_5964 | dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_499 = 6'h37 == replace_index & tag_compare_valid_1 | dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6568 = 6'h38 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_500 = 6'h38 == replace_index & _GEN_5964 | dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_501 = 6'h38 == replace_index & tag_compare_valid_1 | dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6573 = 6'h39 == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_502 = 6'h39 == replace_index & _GEN_5964 | dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_503 = 6'h39 == replace_index & tag_compare_valid_1 | dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6578 = 6'h3a == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_504 = 6'h3a == replace_index & _GEN_5964 | dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_505 = 6'h3a == replace_index & tag_compare_valid_1 | dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6583 = 6'h3b == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_506 = 6'h3b == replace_index & _GEN_5964 | dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_507 = 6'h3b == replace_index & tag_compare_valid_1 | dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6588 = 6'h3c == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_508 = 6'h3c == replace_index & _GEN_5964 | dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_509 = 6'h3c == replace_index & tag_compare_valid_1 | dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6593 = 6'h3d == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_510 = 6'h3d == replace_index & _GEN_5964 | dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_511 = 6'h3d == replace_index & tag_compare_valid_1 | dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6598 = 6'h3e == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_512 = 6'h3e == replace_index & _GEN_5964 | dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_513 = 6'h3e == replace_index & tag_compare_valid_1 | dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_6603 = 6'h3f == replace_index; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_514 = 6'h3f == replace_index & _GEN_5964 | dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_515 = 6'h3f == replace_index & tag_compare_valid_1 | dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 354:{50,50}]
  wire  _GEN_516 = _mmio_read_stall_T ? _GEN_388 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_517 = _mmio_read_stall_T ? _GEN_389 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_518 = _mmio_read_stall_T ? _GEN_390 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_519 = _mmio_read_stall_T ? _GEN_391 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_520 = _mmio_read_stall_T ? _GEN_392 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_521 = _mmio_read_stall_T ? _GEN_393 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_522 = _mmio_read_stall_T ? _GEN_394 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_523 = _mmio_read_stall_T ? _GEN_395 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_524 = _mmio_read_stall_T ? _GEN_396 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_525 = _mmio_read_stall_T ? _GEN_397 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_526 = _mmio_read_stall_T ? _GEN_398 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_527 = _mmio_read_stall_T ? _GEN_399 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_528 = _mmio_read_stall_T ? _GEN_400 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_529 = _mmio_read_stall_T ? _GEN_401 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_530 = _mmio_read_stall_T ? _GEN_402 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_531 = _mmio_read_stall_T ? _GEN_403 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_532 = _mmio_read_stall_T ? _GEN_404 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_533 = _mmio_read_stall_T ? _GEN_405 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_534 = _mmio_read_stall_T ? _GEN_406 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_535 = _mmio_read_stall_T ? _GEN_407 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_536 = _mmio_read_stall_T ? _GEN_408 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_537 = _mmio_read_stall_T ? _GEN_409 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_538 = _mmio_read_stall_T ? _GEN_410 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_539 = _mmio_read_stall_T ? _GEN_411 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_540 = _mmio_read_stall_T ? _GEN_412 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_541 = _mmio_read_stall_T ? _GEN_413 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_542 = _mmio_read_stall_T ? _GEN_414 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_543 = _mmio_read_stall_T ? _GEN_415 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_544 = _mmio_read_stall_T ? _GEN_416 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_545 = _mmio_read_stall_T ? _GEN_417 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_546 = _mmio_read_stall_T ? _GEN_418 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_547 = _mmio_read_stall_T ? _GEN_419 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_548 = _mmio_read_stall_T ? _GEN_420 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_549 = _mmio_read_stall_T ? _GEN_421 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_550 = _mmio_read_stall_T ? _GEN_422 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_551 = _mmio_read_stall_T ? _GEN_423 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_552 = _mmio_read_stall_T ? _GEN_424 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_553 = _mmio_read_stall_T ? _GEN_425 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_554 = _mmio_read_stall_T ? _GEN_426 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_555 = _mmio_read_stall_T ? _GEN_427 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_556 = _mmio_read_stall_T ? _GEN_428 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_557 = _mmio_read_stall_T ? _GEN_429 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_558 = _mmio_read_stall_T ? _GEN_430 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_559 = _mmio_read_stall_T ? _GEN_431 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_560 = _mmio_read_stall_T ? _GEN_432 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_561 = _mmio_read_stall_T ? _GEN_433 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_562 = _mmio_read_stall_T ? _GEN_434 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_563 = _mmio_read_stall_T ? _GEN_435 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_564 = _mmio_read_stall_T ? _GEN_436 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_565 = _mmio_read_stall_T ? _GEN_437 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_566 = _mmio_read_stall_T ? _GEN_438 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_567 = _mmio_read_stall_T ? _GEN_439 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_568 = _mmio_read_stall_T ? _GEN_440 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_569 = _mmio_read_stall_T ? _GEN_441 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_570 = _mmio_read_stall_T ? _GEN_442 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_571 = _mmio_read_stall_T ? _GEN_443 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_572 = _mmio_read_stall_T ? _GEN_444 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_573 = _mmio_read_stall_T ? _GEN_445 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_574 = _mmio_read_stall_T ? _GEN_446 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_575 = _mmio_read_stall_T ? _GEN_447 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_576 = _mmio_read_stall_T ? _GEN_448 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_577 = _mmio_read_stall_T ? _GEN_449 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_578 = _mmio_read_stall_T ? _GEN_450 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_579 = _mmio_read_stall_T ? _GEN_451 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_580 = _mmio_read_stall_T ? _GEN_452 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_581 = _mmio_read_stall_T ? _GEN_453 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_582 = _mmio_read_stall_T ? _GEN_454 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_583 = _mmio_read_stall_T ? _GEN_455 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_584 = _mmio_read_stall_T ? _GEN_456 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_585 = _mmio_read_stall_T ? _GEN_457 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_586 = _mmio_read_stall_T ? _GEN_458 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_587 = _mmio_read_stall_T ? _GEN_459 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_588 = _mmio_read_stall_T ? _GEN_460 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_589 = _mmio_read_stall_T ? _GEN_461 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_590 = _mmio_read_stall_T ? _GEN_462 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_591 = _mmio_read_stall_T ? _GEN_463 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_592 = _mmio_read_stall_T ? _GEN_464 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_593 = _mmio_read_stall_T ? _GEN_465 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_594 = _mmio_read_stall_T ? _GEN_466 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_595 = _mmio_read_stall_T ? _GEN_467 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_596 = _mmio_read_stall_T ? _GEN_468 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_597 = _mmio_read_stall_T ? _GEN_469 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_598 = _mmio_read_stall_T ? _GEN_470 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_599 = _mmio_read_stall_T ? _GEN_471 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_600 = _mmio_read_stall_T ? _GEN_472 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_601 = _mmio_read_stall_T ? _GEN_473 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_602 = _mmio_read_stall_T ? _GEN_474 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_603 = _mmio_read_stall_T ? _GEN_475 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_604 = _mmio_read_stall_T ? _GEN_476 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_605 = _mmio_read_stall_T ? _GEN_477 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_606 = _mmio_read_stall_T ? _GEN_478 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_607 = _mmio_read_stall_T ? _GEN_479 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_608 = _mmio_read_stall_T ? _GEN_480 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_609 = _mmio_read_stall_T ? _GEN_481 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_610 = _mmio_read_stall_T ? _GEN_482 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_611 = _mmio_read_stall_T ? _GEN_483 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_612 = _mmio_read_stall_T ? _GEN_484 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_613 = _mmio_read_stall_T ? _GEN_485 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_614 = _mmio_read_stall_T ? _GEN_486 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_615 = _mmio_read_stall_T ? _GEN_487 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_616 = _mmio_read_stall_T ? _GEN_488 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_617 = _mmio_read_stall_T ? _GEN_489 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_618 = _mmio_read_stall_T ? _GEN_490 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_619 = _mmio_read_stall_T ? _GEN_491 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_620 = _mmio_read_stall_T ? _GEN_492 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_621 = _mmio_read_stall_T ? _GEN_493 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_622 = _mmio_read_stall_T ? _GEN_494 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_623 = _mmio_read_stall_T ? _GEN_495 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_624 = _mmio_read_stall_T ? _GEN_496 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_625 = _mmio_read_stall_T ? _GEN_497 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_626 = _mmio_read_stall_T ? _GEN_498 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_627 = _mmio_read_stall_T ? _GEN_499 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_628 = _mmio_read_stall_T ? _GEN_500 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_629 = _mmio_read_stall_T ? _GEN_501 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_630 = _mmio_read_stall_T ? _GEN_502 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_631 = _mmio_read_stall_T ? _GEN_503 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_632 = _mmio_read_stall_T ? _GEN_504 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_633 = _mmio_read_stall_T ? _GEN_505 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_634 = _mmio_read_stall_T ? _GEN_506 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_635 = _mmio_read_stall_T ? _GEN_507 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_636 = _mmio_read_stall_T ? _GEN_508 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_637 = _mmio_read_stall_T ? _GEN_509 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_638 = _mmio_read_stall_T ? _GEN_510 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_639 = _mmio_read_stall_T ? _GEN_511 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_640 = _mmio_read_stall_T ? _GEN_512 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_641 = _mmio_read_stall_T ? _GEN_513 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_642 = _mmio_read_stall_T ? _GEN_514 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire  _GEN_643 = _mmio_read_stall_T ? _GEN_515 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 353:36]
  wire [63:0] _GEN_644 = _T_7 ? _GEN_15 : saved_rdata; // @[playground/src/cache/DCache.scala 209:28 356:53 357:29]
  wire  _GEN_646 = _io_cpu_dcache_ready_T ? _GEN_324 : lru_0; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_647 = _io_cpu_dcache_ready_T ? _GEN_325 : lru_1; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_648 = _io_cpu_dcache_ready_T ? _GEN_326 : lru_2; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_649 = _io_cpu_dcache_ready_T ? _GEN_327 : lru_3; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_650 = _io_cpu_dcache_ready_T ? _GEN_328 : lru_4; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_651 = _io_cpu_dcache_ready_T ? _GEN_329 : lru_5; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_652 = _io_cpu_dcache_ready_T ? _GEN_330 : lru_6; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_653 = _io_cpu_dcache_ready_T ? _GEN_331 : lru_7; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_654 = _io_cpu_dcache_ready_T ? _GEN_332 : lru_8; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_655 = _io_cpu_dcache_ready_T ? _GEN_333 : lru_9; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_656 = _io_cpu_dcache_ready_T ? _GEN_334 : lru_10; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_657 = _io_cpu_dcache_ready_T ? _GEN_335 : lru_11; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_658 = _io_cpu_dcache_ready_T ? _GEN_336 : lru_12; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_659 = _io_cpu_dcache_ready_T ? _GEN_337 : lru_13; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_660 = _io_cpu_dcache_ready_T ? _GEN_338 : lru_14; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_661 = _io_cpu_dcache_ready_T ? _GEN_339 : lru_15; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_662 = _io_cpu_dcache_ready_T ? _GEN_340 : lru_16; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_663 = _io_cpu_dcache_ready_T ? _GEN_341 : lru_17; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_664 = _io_cpu_dcache_ready_T ? _GEN_342 : lru_18; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_665 = _io_cpu_dcache_ready_T ? _GEN_343 : lru_19; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_666 = _io_cpu_dcache_ready_T ? _GEN_344 : lru_20; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_667 = _io_cpu_dcache_ready_T ? _GEN_345 : lru_21; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_668 = _io_cpu_dcache_ready_T ? _GEN_346 : lru_22; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_669 = _io_cpu_dcache_ready_T ? _GEN_347 : lru_23; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_670 = _io_cpu_dcache_ready_T ? _GEN_348 : lru_24; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_671 = _io_cpu_dcache_ready_T ? _GEN_349 : lru_25; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_672 = _io_cpu_dcache_ready_T ? _GEN_350 : lru_26; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_673 = _io_cpu_dcache_ready_T ? _GEN_351 : lru_27; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_674 = _io_cpu_dcache_ready_T ? _GEN_352 : lru_28; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_675 = _io_cpu_dcache_ready_T ? _GEN_353 : lru_29; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_676 = _io_cpu_dcache_ready_T ? _GEN_354 : lru_30; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_677 = _io_cpu_dcache_ready_T ? _GEN_355 : lru_31; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_678 = _io_cpu_dcache_ready_T ? _GEN_356 : lru_32; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_679 = _io_cpu_dcache_ready_T ? _GEN_357 : lru_33; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_680 = _io_cpu_dcache_ready_T ? _GEN_358 : lru_34; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_681 = _io_cpu_dcache_ready_T ? _GEN_359 : lru_35; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_682 = _io_cpu_dcache_ready_T ? _GEN_360 : lru_36; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_683 = _io_cpu_dcache_ready_T ? _GEN_361 : lru_37; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_684 = _io_cpu_dcache_ready_T ? _GEN_362 : lru_38; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_685 = _io_cpu_dcache_ready_T ? _GEN_363 : lru_39; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_686 = _io_cpu_dcache_ready_T ? _GEN_364 : lru_40; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_687 = _io_cpu_dcache_ready_T ? _GEN_365 : lru_41; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_688 = _io_cpu_dcache_ready_T ? _GEN_366 : lru_42; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_689 = _io_cpu_dcache_ready_T ? _GEN_367 : lru_43; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_690 = _io_cpu_dcache_ready_T ? _GEN_368 : lru_44; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_691 = _io_cpu_dcache_ready_T ? _GEN_369 : lru_45; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_692 = _io_cpu_dcache_ready_T ? _GEN_370 : lru_46; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_693 = _io_cpu_dcache_ready_T ? _GEN_371 : lru_47; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_694 = _io_cpu_dcache_ready_T ? _GEN_372 : lru_48; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_695 = _io_cpu_dcache_ready_T ? _GEN_373 : lru_49; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_696 = _io_cpu_dcache_ready_T ? _GEN_374 : lru_50; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_697 = _io_cpu_dcache_ready_T ? _GEN_375 : lru_51; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_698 = _io_cpu_dcache_ready_T ? _GEN_376 : lru_52; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_699 = _io_cpu_dcache_ready_T ? _GEN_377 : lru_53; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_700 = _io_cpu_dcache_ready_T ? _GEN_378 : lru_54; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_701 = _io_cpu_dcache_ready_T ? _GEN_379 : lru_55; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_702 = _io_cpu_dcache_ready_T ? _GEN_380 : lru_56; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_703 = _io_cpu_dcache_ready_T ? _GEN_381 : lru_57; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_704 = _io_cpu_dcache_ready_T ? _GEN_382 : lru_58; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_705 = _io_cpu_dcache_ready_T ? _GEN_383 : lru_59; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_706 = _io_cpu_dcache_ready_T ? _GEN_384 : lru_60; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_707 = _io_cpu_dcache_ready_T ? _GEN_385 : lru_61; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_708 = _io_cpu_dcache_ready_T ? _GEN_386 : lru_62; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_709 = _io_cpu_dcache_ready_T ? _GEN_387 : lru_63; // @[playground/src/cache/DCache.scala 136:22 350:33]
  wire  _GEN_710 = _io_cpu_dcache_ready_T ? _GEN_516 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_711 = _io_cpu_dcache_ready_T ? _GEN_517 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_712 = _io_cpu_dcache_ready_T ? _GEN_518 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_713 = _io_cpu_dcache_ready_T ? _GEN_519 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_714 = _io_cpu_dcache_ready_T ? _GEN_520 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_715 = _io_cpu_dcache_ready_T ? _GEN_521 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_716 = _io_cpu_dcache_ready_T ? _GEN_522 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_717 = _io_cpu_dcache_ready_T ? _GEN_523 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_718 = _io_cpu_dcache_ready_T ? _GEN_524 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_719 = _io_cpu_dcache_ready_T ? _GEN_525 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_720 = _io_cpu_dcache_ready_T ? _GEN_526 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_721 = _io_cpu_dcache_ready_T ? _GEN_527 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_722 = _io_cpu_dcache_ready_T ? _GEN_528 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_723 = _io_cpu_dcache_ready_T ? _GEN_529 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_724 = _io_cpu_dcache_ready_T ? _GEN_530 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_725 = _io_cpu_dcache_ready_T ? _GEN_531 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_726 = _io_cpu_dcache_ready_T ? _GEN_532 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_727 = _io_cpu_dcache_ready_T ? _GEN_533 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_728 = _io_cpu_dcache_ready_T ? _GEN_534 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_729 = _io_cpu_dcache_ready_T ? _GEN_535 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_730 = _io_cpu_dcache_ready_T ? _GEN_536 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_731 = _io_cpu_dcache_ready_T ? _GEN_537 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_732 = _io_cpu_dcache_ready_T ? _GEN_538 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_733 = _io_cpu_dcache_ready_T ? _GEN_539 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_734 = _io_cpu_dcache_ready_T ? _GEN_540 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_735 = _io_cpu_dcache_ready_T ? _GEN_541 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_736 = _io_cpu_dcache_ready_T ? _GEN_542 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_737 = _io_cpu_dcache_ready_T ? _GEN_543 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_738 = _io_cpu_dcache_ready_T ? _GEN_544 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_739 = _io_cpu_dcache_ready_T ? _GEN_545 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_740 = _io_cpu_dcache_ready_T ? _GEN_546 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_741 = _io_cpu_dcache_ready_T ? _GEN_547 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_742 = _io_cpu_dcache_ready_T ? _GEN_548 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_743 = _io_cpu_dcache_ready_T ? _GEN_549 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_744 = _io_cpu_dcache_ready_T ? _GEN_550 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_745 = _io_cpu_dcache_ready_T ? _GEN_551 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_746 = _io_cpu_dcache_ready_T ? _GEN_552 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_747 = _io_cpu_dcache_ready_T ? _GEN_553 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_748 = _io_cpu_dcache_ready_T ? _GEN_554 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_749 = _io_cpu_dcache_ready_T ? _GEN_555 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_750 = _io_cpu_dcache_ready_T ? _GEN_556 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_751 = _io_cpu_dcache_ready_T ? _GEN_557 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_752 = _io_cpu_dcache_ready_T ? _GEN_558 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_753 = _io_cpu_dcache_ready_T ? _GEN_559 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_754 = _io_cpu_dcache_ready_T ? _GEN_560 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_755 = _io_cpu_dcache_ready_T ? _GEN_561 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_756 = _io_cpu_dcache_ready_T ? _GEN_562 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_757 = _io_cpu_dcache_ready_T ? _GEN_563 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_758 = _io_cpu_dcache_ready_T ? _GEN_564 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_759 = _io_cpu_dcache_ready_T ? _GEN_565 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_760 = _io_cpu_dcache_ready_T ? _GEN_566 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_761 = _io_cpu_dcache_ready_T ? _GEN_567 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_762 = _io_cpu_dcache_ready_T ? _GEN_568 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_763 = _io_cpu_dcache_ready_T ? _GEN_569 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_764 = _io_cpu_dcache_ready_T ? _GEN_570 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_765 = _io_cpu_dcache_ready_T ? _GEN_571 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_766 = _io_cpu_dcache_ready_T ? _GEN_572 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_767 = _io_cpu_dcache_ready_T ? _GEN_573 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_768 = _io_cpu_dcache_ready_T ? _GEN_574 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_769 = _io_cpu_dcache_ready_T ? _GEN_575 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_770 = _io_cpu_dcache_ready_T ? _GEN_576 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_771 = _io_cpu_dcache_ready_T ? _GEN_577 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_772 = _io_cpu_dcache_ready_T ? _GEN_578 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_773 = _io_cpu_dcache_ready_T ? _GEN_579 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_774 = _io_cpu_dcache_ready_T ? _GEN_580 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_775 = _io_cpu_dcache_ready_T ? _GEN_581 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_776 = _io_cpu_dcache_ready_T ? _GEN_582 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_777 = _io_cpu_dcache_ready_T ? _GEN_583 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_778 = _io_cpu_dcache_ready_T ? _GEN_584 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_779 = _io_cpu_dcache_ready_T ? _GEN_585 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_780 = _io_cpu_dcache_ready_T ? _GEN_586 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_781 = _io_cpu_dcache_ready_T ? _GEN_587 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_782 = _io_cpu_dcache_ready_T ? _GEN_588 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_783 = _io_cpu_dcache_ready_T ? _GEN_589 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_784 = _io_cpu_dcache_ready_T ? _GEN_590 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_785 = _io_cpu_dcache_ready_T ? _GEN_591 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_786 = _io_cpu_dcache_ready_T ? _GEN_592 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_787 = _io_cpu_dcache_ready_T ? _GEN_593 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_788 = _io_cpu_dcache_ready_T ? _GEN_594 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_789 = _io_cpu_dcache_ready_T ? _GEN_595 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_790 = _io_cpu_dcache_ready_T ? _GEN_596 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_791 = _io_cpu_dcache_ready_T ? _GEN_597 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_792 = _io_cpu_dcache_ready_T ? _GEN_598 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_793 = _io_cpu_dcache_ready_T ? _GEN_599 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_794 = _io_cpu_dcache_ready_T ? _GEN_600 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_795 = _io_cpu_dcache_ready_T ? _GEN_601 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_796 = _io_cpu_dcache_ready_T ? _GEN_602 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_797 = _io_cpu_dcache_ready_T ? _GEN_603 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_798 = _io_cpu_dcache_ready_T ? _GEN_604 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_799 = _io_cpu_dcache_ready_T ? _GEN_605 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_800 = _io_cpu_dcache_ready_T ? _GEN_606 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_801 = _io_cpu_dcache_ready_T ? _GEN_607 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_802 = _io_cpu_dcache_ready_T ? _GEN_608 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_803 = _io_cpu_dcache_ready_T ? _GEN_609 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_804 = _io_cpu_dcache_ready_T ? _GEN_610 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_805 = _io_cpu_dcache_ready_T ? _GEN_611 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_806 = _io_cpu_dcache_ready_T ? _GEN_612 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_807 = _io_cpu_dcache_ready_T ? _GEN_613 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_808 = _io_cpu_dcache_ready_T ? _GEN_614 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_809 = _io_cpu_dcache_ready_T ? _GEN_615 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_810 = _io_cpu_dcache_ready_T ? _GEN_616 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_811 = _io_cpu_dcache_ready_T ? _GEN_617 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_812 = _io_cpu_dcache_ready_T ? _GEN_618 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_813 = _io_cpu_dcache_ready_T ? _GEN_619 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_814 = _io_cpu_dcache_ready_T ? _GEN_620 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_815 = _io_cpu_dcache_ready_T ? _GEN_621 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_816 = _io_cpu_dcache_ready_T ? _GEN_622 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_817 = _io_cpu_dcache_ready_T ? _GEN_623 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_818 = _io_cpu_dcache_ready_T ? _GEN_624 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_819 = _io_cpu_dcache_ready_T ? _GEN_625 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_820 = _io_cpu_dcache_ready_T ? _GEN_626 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_821 = _io_cpu_dcache_ready_T ? _GEN_627 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_822 = _io_cpu_dcache_ready_T ? _GEN_628 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_823 = _io_cpu_dcache_ready_T ? _GEN_629 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_824 = _io_cpu_dcache_ready_T ? _GEN_630 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_825 = _io_cpu_dcache_ready_T ? _GEN_631 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_826 = _io_cpu_dcache_ready_T ? _GEN_632 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_827 = _io_cpu_dcache_ready_T ? _GEN_633 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_828 = _io_cpu_dcache_ready_T ? _GEN_634 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_829 = _io_cpu_dcache_ready_T ? _GEN_635 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_830 = _io_cpu_dcache_ready_T ? _GEN_636 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_831 = _io_cpu_dcache_ready_T ? _GEN_637 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_832 = _io_cpu_dcache_ready_T ? _GEN_638 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_833 = _io_cpu_dcache_ready_T ? _GEN_639 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_834 = _io_cpu_dcache_ready_T ? _GEN_640 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_835 = _io_cpu_dcache_ready_T ? _GEN_641 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_836 = _io_cpu_dcache_ready_T ? _GEN_642 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire  _GEN_837 = _io_cpu_dcache_ready_T ? _GEN_643 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 350:33]
  wire [63:0] _GEN_838 = _io_cpu_dcache_ready_T ? _GEN_644 : saved_rdata; // @[playground/src/cache/DCache.scala 209:28 350:33]
  wire [2:0] _GEN_839 = _io_cpu_dcache_ready_T ? _GEN_300 : state; // @[playground/src/cache/DCache.scala 350:33 90:94]
  wire [2:0] _GEN_840 = _cached_stall_T_1 ? 3'h3 : _GEN_839; // @[playground/src/cache/DCache.scala 347:28 348:19]
  wire  _GEN_841 = _cached_stall_T_1 ? lru_0 : _GEN_646; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_842 = _cached_stall_T_1 ? lru_1 : _GEN_647; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_843 = _cached_stall_T_1 ? lru_2 : _GEN_648; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_844 = _cached_stall_T_1 ? lru_3 : _GEN_649; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_845 = _cached_stall_T_1 ? lru_4 : _GEN_650; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_846 = _cached_stall_T_1 ? lru_5 : _GEN_651; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_847 = _cached_stall_T_1 ? lru_6 : _GEN_652; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_848 = _cached_stall_T_1 ? lru_7 : _GEN_653; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_849 = _cached_stall_T_1 ? lru_8 : _GEN_654; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_850 = _cached_stall_T_1 ? lru_9 : _GEN_655; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_851 = _cached_stall_T_1 ? lru_10 : _GEN_656; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_852 = _cached_stall_T_1 ? lru_11 : _GEN_657; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_853 = _cached_stall_T_1 ? lru_12 : _GEN_658; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_854 = _cached_stall_T_1 ? lru_13 : _GEN_659; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_855 = _cached_stall_T_1 ? lru_14 : _GEN_660; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_856 = _cached_stall_T_1 ? lru_15 : _GEN_661; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_857 = _cached_stall_T_1 ? lru_16 : _GEN_662; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_858 = _cached_stall_T_1 ? lru_17 : _GEN_663; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_859 = _cached_stall_T_1 ? lru_18 : _GEN_664; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_860 = _cached_stall_T_1 ? lru_19 : _GEN_665; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_861 = _cached_stall_T_1 ? lru_20 : _GEN_666; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_862 = _cached_stall_T_1 ? lru_21 : _GEN_667; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_863 = _cached_stall_T_1 ? lru_22 : _GEN_668; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_864 = _cached_stall_T_1 ? lru_23 : _GEN_669; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_865 = _cached_stall_T_1 ? lru_24 : _GEN_670; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_866 = _cached_stall_T_1 ? lru_25 : _GEN_671; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_867 = _cached_stall_T_1 ? lru_26 : _GEN_672; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_868 = _cached_stall_T_1 ? lru_27 : _GEN_673; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_869 = _cached_stall_T_1 ? lru_28 : _GEN_674; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_870 = _cached_stall_T_1 ? lru_29 : _GEN_675; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_871 = _cached_stall_T_1 ? lru_30 : _GEN_676; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_872 = _cached_stall_T_1 ? lru_31 : _GEN_677; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_873 = _cached_stall_T_1 ? lru_32 : _GEN_678; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_874 = _cached_stall_T_1 ? lru_33 : _GEN_679; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_875 = _cached_stall_T_1 ? lru_34 : _GEN_680; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_876 = _cached_stall_T_1 ? lru_35 : _GEN_681; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_877 = _cached_stall_T_1 ? lru_36 : _GEN_682; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_878 = _cached_stall_T_1 ? lru_37 : _GEN_683; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_879 = _cached_stall_T_1 ? lru_38 : _GEN_684; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_880 = _cached_stall_T_1 ? lru_39 : _GEN_685; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_881 = _cached_stall_T_1 ? lru_40 : _GEN_686; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_882 = _cached_stall_T_1 ? lru_41 : _GEN_687; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_883 = _cached_stall_T_1 ? lru_42 : _GEN_688; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_884 = _cached_stall_T_1 ? lru_43 : _GEN_689; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_885 = _cached_stall_T_1 ? lru_44 : _GEN_690; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_886 = _cached_stall_T_1 ? lru_45 : _GEN_691; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_887 = _cached_stall_T_1 ? lru_46 : _GEN_692; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_888 = _cached_stall_T_1 ? lru_47 : _GEN_693; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_889 = _cached_stall_T_1 ? lru_48 : _GEN_694; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_890 = _cached_stall_T_1 ? lru_49 : _GEN_695; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_891 = _cached_stall_T_1 ? lru_50 : _GEN_696; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_892 = _cached_stall_T_1 ? lru_51 : _GEN_697; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_893 = _cached_stall_T_1 ? lru_52 : _GEN_698; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_894 = _cached_stall_T_1 ? lru_53 : _GEN_699; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_895 = _cached_stall_T_1 ? lru_54 : _GEN_700; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_896 = _cached_stall_T_1 ? lru_55 : _GEN_701; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_897 = _cached_stall_T_1 ? lru_56 : _GEN_702; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_898 = _cached_stall_T_1 ? lru_57 : _GEN_703; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_899 = _cached_stall_T_1 ? lru_58 : _GEN_704; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_900 = _cached_stall_T_1 ? lru_59 : _GEN_705; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_901 = _cached_stall_T_1 ? lru_60 : _GEN_706; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_902 = _cached_stall_T_1 ? lru_61 : _GEN_707; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_903 = _cached_stall_T_1 ? lru_62 : _GEN_708; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_904 = _cached_stall_T_1 ? lru_63 : _GEN_709; // @[playground/src/cache/DCache.scala 136:22 347:28]
  wire  _GEN_905 = _cached_stall_T_1 ? dirty_0_0 : _GEN_710; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_906 = _cached_stall_T_1 ? dirty_0_1 : _GEN_711; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_907 = _cached_stall_T_1 ? dirty_1_0 : _GEN_712; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_908 = _cached_stall_T_1 ? dirty_1_1 : _GEN_713; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_909 = _cached_stall_T_1 ? dirty_2_0 : _GEN_714; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_910 = _cached_stall_T_1 ? dirty_2_1 : _GEN_715; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_911 = _cached_stall_T_1 ? dirty_3_0 : _GEN_716; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_912 = _cached_stall_T_1 ? dirty_3_1 : _GEN_717; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_913 = _cached_stall_T_1 ? dirty_4_0 : _GEN_718; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_914 = _cached_stall_T_1 ? dirty_4_1 : _GEN_719; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_915 = _cached_stall_T_1 ? dirty_5_0 : _GEN_720; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_916 = _cached_stall_T_1 ? dirty_5_1 : _GEN_721; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_917 = _cached_stall_T_1 ? dirty_6_0 : _GEN_722; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_918 = _cached_stall_T_1 ? dirty_6_1 : _GEN_723; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_919 = _cached_stall_T_1 ? dirty_7_0 : _GEN_724; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_920 = _cached_stall_T_1 ? dirty_7_1 : _GEN_725; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_921 = _cached_stall_T_1 ? dirty_8_0 : _GEN_726; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_922 = _cached_stall_T_1 ? dirty_8_1 : _GEN_727; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_923 = _cached_stall_T_1 ? dirty_9_0 : _GEN_728; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_924 = _cached_stall_T_1 ? dirty_9_1 : _GEN_729; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_925 = _cached_stall_T_1 ? dirty_10_0 : _GEN_730; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_926 = _cached_stall_T_1 ? dirty_10_1 : _GEN_731; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_927 = _cached_stall_T_1 ? dirty_11_0 : _GEN_732; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_928 = _cached_stall_T_1 ? dirty_11_1 : _GEN_733; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_929 = _cached_stall_T_1 ? dirty_12_0 : _GEN_734; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_930 = _cached_stall_T_1 ? dirty_12_1 : _GEN_735; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_931 = _cached_stall_T_1 ? dirty_13_0 : _GEN_736; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_932 = _cached_stall_T_1 ? dirty_13_1 : _GEN_737; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_933 = _cached_stall_T_1 ? dirty_14_0 : _GEN_738; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_934 = _cached_stall_T_1 ? dirty_14_1 : _GEN_739; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_935 = _cached_stall_T_1 ? dirty_15_0 : _GEN_740; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_936 = _cached_stall_T_1 ? dirty_15_1 : _GEN_741; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_937 = _cached_stall_T_1 ? dirty_16_0 : _GEN_742; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_938 = _cached_stall_T_1 ? dirty_16_1 : _GEN_743; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_939 = _cached_stall_T_1 ? dirty_17_0 : _GEN_744; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_940 = _cached_stall_T_1 ? dirty_17_1 : _GEN_745; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_941 = _cached_stall_T_1 ? dirty_18_0 : _GEN_746; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_942 = _cached_stall_T_1 ? dirty_18_1 : _GEN_747; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_943 = _cached_stall_T_1 ? dirty_19_0 : _GEN_748; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_944 = _cached_stall_T_1 ? dirty_19_1 : _GEN_749; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_945 = _cached_stall_T_1 ? dirty_20_0 : _GEN_750; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_946 = _cached_stall_T_1 ? dirty_20_1 : _GEN_751; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_947 = _cached_stall_T_1 ? dirty_21_0 : _GEN_752; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_948 = _cached_stall_T_1 ? dirty_21_1 : _GEN_753; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_949 = _cached_stall_T_1 ? dirty_22_0 : _GEN_754; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_950 = _cached_stall_T_1 ? dirty_22_1 : _GEN_755; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_951 = _cached_stall_T_1 ? dirty_23_0 : _GEN_756; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_952 = _cached_stall_T_1 ? dirty_23_1 : _GEN_757; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_953 = _cached_stall_T_1 ? dirty_24_0 : _GEN_758; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_954 = _cached_stall_T_1 ? dirty_24_1 : _GEN_759; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_955 = _cached_stall_T_1 ? dirty_25_0 : _GEN_760; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_956 = _cached_stall_T_1 ? dirty_25_1 : _GEN_761; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_957 = _cached_stall_T_1 ? dirty_26_0 : _GEN_762; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_958 = _cached_stall_T_1 ? dirty_26_1 : _GEN_763; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_959 = _cached_stall_T_1 ? dirty_27_0 : _GEN_764; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_960 = _cached_stall_T_1 ? dirty_27_1 : _GEN_765; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_961 = _cached_stall_T_1 ? dirty_28_0 : _GEN_766; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_962 = _cached_stall_T_1 ? dirty_28_1 : _GEN_767; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_963 = _cached_stall_T_1 ? dirty_29_0 : _GEN_768; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_964 = _cached_stall_T_1 ? dirty_29_1 : _GEN_769; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_965 = _cached_stall_T_1 ? dirty_30_0 : _GEN_770; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_966 = _cached_stall_T_1 ? dirty_30_1 : _GEN_771; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_967 = _cached_stall_T_1 ? dirty_31_0 : _GEN_772; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_968 = _cached_stall_T_1 ? dirty_31_1 : _GEN_773; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_969 = _cached_stall_T_1 ? dirty_32_0 : _GEN_774; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_970 = _cached_stall_T_1 ? dirty_32_1 : _GEN_775; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_971 = _cached_stall_T_1 ? dirty_33_0 : _GEN_776; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_972 = _cached_stall_T_1 ? dirty_33_1 : _GEN_777; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_973 = _cached_stall_T_1 ? dirty_34_0 : _GEN_778; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_974 = _cached_stall_T_1 ? dirty_34_1 : _GEN_779; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_975 = _cached_stall_T_1 ? dirty_35_0 : _GEN_780; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_976 = _cached_stall_T_1 ? dirty_35_1 : _GEN_781; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_977 = _cached_stall_T_1 ? dirty_36_0 : _GEN_782; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_978 = _cached_stall_T_1 ? dirty_36_1 : _GEN_783; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_979 = _cached_stall_T_1 ? dirty_37_0 : _GEN_784; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_980 = _cached_stall_T_1 ? dirty_37_1 : _GEN_785; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_981 = _cached_stall_T_1 ? dirty_38_0 : _GEN_786; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_982 = _cached_stall_T_1 ? dirty_38_1 : _GEN_787; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_983 = _cached_stall_T_1 ? dirty_39_0 : _GEN_788; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_984 = _cached_stall_T_1 ? dirty_39_1 : _GEN_789; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_985 = _cached_stall_T_1 ? dirty_40_0 : _GEN_790; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_986 = _cached_stall_T_1 ? dirty_40_1 : _GEN_791; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_987 = _cached_stall_T_1 ? dirty_41_0 : _GEN_792; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_988 = _cached_stall_T_1 ? dirty_41_1 : _GEN_793; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_989 = _cached_stall_T_1 ? dirty_42_0 : _GEN_794; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_990 = _cached_stall_T_1 ? dirty_42_1 : _GEN_795; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_991 = _cached_stall_T_1 ? dirty_43_0 : _GEN_796; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_992 = _cached_stall_T_1 ? dirty_43_1 : _GEN_797; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_993 = _cached_stall_T_1 ? dirty_44_0 : _GEN_798; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_994 = _cached_stall_T_1 ? dirty_44_1 : _GEN_799; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_995 = _cached_stall_T_1 ? dirty_45_0 : _GEN_800; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_996 = _cached_stall_T_1 ? dirty_45_1 : _GEN_801; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_997 = _cached_stall_T_1 ? dirty_46_0 : _GEN_802; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_998 = _cached_stall_T_1 ? dirty_46_1 : _GEN_803; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_999 = _cached_stall_T_1 ? dirty_47_0 : _GEN_804; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1000 = _cached_stall_T_1 ? dirty_47_1 : _GEN_805; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1001 = _cached_stall_T_1 ? dirty_48_0 : _GEN_806; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1002 = _cached_stall_T_1 ? dirty_48_1 : _GEN_807; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1003 = _cached_stall_T_1 ? dirty_49_0 : _GEN_808; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1004 = _cached_stall_T_1 ? dirty_49_1 : _GEN_809; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1005 = _cached_stall_T_1 ? dirty_50_0 : _GEN_810; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1006 = _cached_stall_T_1 ? dirty_50_1 : _GEN_811; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1007 = _cached_stall_T_1 ? dirty_51_0 : _GEN_812; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1008 = _cached_stall_T_1 ? dirty_51_1 : _GEN_813; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1009 = _cached_stall_T_1 ? dirty_52_0 : _GEN_814; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1010 = _cached_stall_T_1 ? dirty_52_1 : _GEN_815; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1011 = _cached_stall_T_1 ? dirty_53_0 : _GEN_816; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1012 = _cached_stall_T_1 ? dirty_53_1 : _GEN_817; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1013 = _cached_stall_T_1 ? dirty_54_0 : _GEN_818; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1014 = _cached_stall_T_1 ? dirty_54_1 : _GEN_819; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1015 = _cached_stall_T_1 ? dirty_55_0 : _GEN_820; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1016 = _cached_stall_T_1 ? dirty_55_1 : _GEN_821; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1017 = _cached_stall_T_1 ? dirty_56_0 : _GEN_822; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1018 = _cached_stall_T_1 ? dirty_56_1 : _GEN_823; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1019 = _cached_stall_T_1 ? dirty_57_0 : _GEN_824; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1020 = _cached_stall_T_1 ? dirty_57_1 : _GEN_825; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1021 = _cached_stall_T_1 ? dirty_58_0 : _GEN_826; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1022 = _cached_stall_T_1 ? dirty_58_1 : _GEN_827; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1023 = _cached_stall_T_1 ? dirty_59_0 : _GEN_828; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1024 = _cached_stall_T_1 ? dirty_59_1 : _GEN_829; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1025 = _cached_stall_T_1 ? dirty_60_0 : _GEN_830; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1026 = _cached_stall_T_1 ? dirty_60_1 : _GEN_831; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1027 = _cached_stall_T_1 ? dirty_61_0 : _GEN_832; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1028 = _cached_stall_T_1 ? dirty_61_1 : _GEN_833; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1029 = _cached_stall_T_1 ? dirty_62_0 : _GEN_834; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1030 = _cached_stall_T_1 ? dirty_62_1 : _GEN_835; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1031 = _cached_stall_T_1 ? dirty_63_0 : _GEN_836; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire  _GEN_1032 = _cached_stall_T_1 ? dirty_63_1 : _GEN_837; // @[playground/src/cache/DCache.scala 135:22 347:28]
  wire [63:0] _GEN_1033 = _cached_stall_T_1 ? saved_rdata : _GEN_838; // @[playground/src/cache/DCache.scala 209:28 347:28]
  wire  _GEN_1034 = io_cpu_tlb_uncached & _GEN_313; // @[playground/src/cache/DCache.scala 155:26 325:41]
  wire [63:0] _GEN_1035 = io_cpu_tlb_uncached ? _GEN_314 : 64'h0; // @[playground/src/cache/DCache.scala 156:26 325:41]
  wire [7:0] _GEN_1036 = io_cpu_tlb_uncached ? _GEN_315 : 8'h0; // @[playground/src/cache/DCache.scala 156:26 325:41]
  wire [7:0] _GEN_1037 = io_cpu_tlb_uncached ? _GEN_316 : 8'h0; // @[playground/src/cache/DCache.scala 156:26 325:41]
  wire [63:0] _GEN_1038 = io_cpu_tlb_uncached ? _GEN_317 : 64'h0; // @[playground/src/cache/DCache.scala 156:26 325:41]
  wire [2:0] _GEN_1039 = io_cpu_tlb_uncached ? _GEN_318 : _GEN_840; // @[playground/src/cache/DCache.scala 325:41]
  wire [31:0] _GEN_1040 = io_cpu_tlb_uncached ? _GEN_319 : ar_addr; // @[playground/src/cache/DCache.scala 259:24 325:41]
  wire [7:0] _GEN_1041 = io_cpu_tlb_uncached ? _GEN_320 : ar_len; // @[playground/src/cache/DCache.scala 259:24 325:41]
  wire [7:0] _GEN_1042 = io_cpu_tlb_uncached ? _GEN_321 : {{5'd0}, ar_size}; // @[playground/src/cache/DCache.scala 259:24 325:41]
  wire  _GEN_1043 = io_cpu_tlb_uncached ? _GEN_322 : arvalid; // @[playground/src/cache/DCache.scala 260:24 325:41]
  wire  _GEN_1044 = io_cpu_tlb_uncached ? _GEN_323 : rready; // @[playground/src/cache/DCache.scala 263:23 325:41]
  wire  _GEN_1045 = io_cpu_tlb_uncached ? lru_0 : _GEN_841; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1046 = io_cpu_tlb_uncached ? lru_1 : _GEN_842; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1047 = io_cpu_tlb_uncached ? lru_2 : _GEN_843; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1048 = io_cpu_tlb_uncached ? lru_3 : _GEN_844; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1049 = io_cpu_tlb_uncached ? lru_4 : _GEN_845; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1050 = io_cpu_tlb_uncached ? lru_5 : _GEN_846; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1051 = io_cpu_tlb_uncached ? lru_6 : _GEN_847; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1052 = io_cpu_tlb_uncached ? lru_7 : _GEN_848; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1053 = io_cpu_tlb_uncached ? lru_8 : _GEN_849; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1054 = io_cpu_tlb_uncached ? lru_9 : _GEN_850; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1055 = io_cpu_tlb_uncached ? lru_10 : _GEN_851; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1056 = io_cpu_tlb_uncached ? lru_11 : _GEN_852; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1057 = io_cpu_tlb_uncached ? lru_12 : _GEN_853; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1058 = io_cpu_tlb_uncached ? lru_13 : _GEN_854; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1059 = io_cpu_tlb_uncached ? lru_14 : _GEN_855; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1060 = io_cpu_tlb_uncached ? lru_15 : _GEN_856; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1061 = io_cpu_tlb_uncached ? lru_16 : _GEN_857; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1062 = io_cpu_tlb_uncached ? lru_17 : _GEN_858; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1063 = io_cpu_tlb_uncached ? lru_18 : _GEN_859; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1064 = io_cpu_tlb_uncached ? lru_19 : _GEN_860; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1065 = io_cpu_tlb_uncached ? lru_20 : _GEN_861; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1066 = io_cpu_tlb_uncached ? lru_21 : _GEN_862; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1067 = io_cpu_tlb_uncached ? lru_22 : _GEN_863; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1068 = io_cpu_tlb_uncached ? lru_23 : _GEN_864; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1069 = io_cpu_tlb_uncached ? lru_24 : _GEN_865; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1070 = io_cpu_tlb_uncached ? lru_25 : _GEN_866; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1071 = io_cpu_tlb_uncached ? lru_26 : _GEN_867; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1072 = io_cpu_tlb_uncached ? lru_27 : _GEN_868; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1073 = io_cpu_tlb_uncached ? lru_28 : _GEN_869; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1074 = io_cpu_tlb_uncached ? lru_29 : _GEN_870; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1075 = io_cpu_tlb_uncached ? lru_30 : _GEN_871; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1076 = io_cpu_tlb_uncached ? lru_31 : _GEN_872; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1077 = io_cpu_tlb_uncached ? lru_32 : _GEN_873; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1078 = io_cpu_tlb_uncached ? lru_33 : _GEN_874; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1079 = io_cpu_tlb_uncached ? lru_34 : _GEN_875; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1080 = io_cpu_tlb_uncached ? lru_35 : _GEN_876; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1081 = io_cpu_tlb_uncached ? lru_36 : _GEN_877; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1082 = io_cpu_tlb_uncached ? lru_37 : _GEN_878; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1083 = io_cpu_tlb_uncached ? lru_38 : _GEN_879; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1084 = io_cpu_tlb_uncached ? lru_39 : _GEN_880; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1085 = io_cpu_tlb_uncached ? lru_40 : _GEN_881; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1086 = io_cpu_tlb_uncached ? lru_41 : _GEN_882; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1087 = io_cpu_tlb_uncached ? lru_42 : _GEN_883; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1088 = io_cpu_tlb_uncached ? lru_43 : _GEN_884; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1089 = io_cpu_tlb_uncached ? lru_44 : _GEN_885; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1090 = io_cpu_tlb_uncached ? lru_45 : _GEN_886; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1091 = io_cpu_tlb_uncached ? lru_46 : _GEN_887; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1092 = io_cpu_tlb_uncached ? lru_47 : _GEN_888; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1093 = io_cpu_tlb_uncached ? lru_48 : _GEN_889; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1094 = io_cpu_tlb_uncached ? lru_49 : _GEN_890; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1095 = io_cpu_tlb_uncached ? lru_50 : _GEN_891; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1096 = io_cpu_tlb_uncached ? lru_51 : _GEN_892; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1097 = io_cpu_tlb_uncached ? lru_52 : _GEN_893; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1098 = io_cpu_tlb_uncached ? lru_53 : _GEN_894; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1099 = io_cpu_tlb_uncached ? lru_54 : _GEN_895; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1100 = io_cpu_tlb_uncached ? lru_55 : _GEN_896; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1101 = io_cpu_tlb_uncached ? lru_56 : _GEN_897; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1102 = io_cpu_tlb_uncached ? lru_57 : _GEN_898; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1103 = io_cpu_tlb_uncached ? lru_58 : _GEN_899; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1104 = io_cpu_tlb_uncached ? lru_59 : _GEN_900; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1105 = io_cpu_tlb_uncached ? lru_60 : _GEN_901; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1106 = io_cpu_tlb_uncached ? lru_61 : _GEN_902; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1107 = io_cpu_tlb_uncached ? lru_62 : _GEN_903; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1108 = io_cpu_tlb_uncached ? lru_63 : _GEN_904; // @[playground/src/cache/DCache.scala 136:22 325:41]
  wire  _GEN_1109 = io_cpu_tlb_uncached ? dirty_0_0 : _GEN_905; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1110 = io_cpu_tlb_uncached ? dirty_0_1 : _GEN_906; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1111 = io_cpu_tlb_uncached ? dirty_1_0 : _GEN_907; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1112 = io_cpu_tlb_uncached ? dirty_1_1 : _GEN_908; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1113 = io_cpu_tlb_uncached ? dirty_2_0 : _GEN_909; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1114 = io_cpu_tlb_uncached ? dirty_2_1 : _GEN_910; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1115 = io_cpu_tlb_uncached ? dirty_3_0 : _GEN_911; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1116 = io_cpu_tlb_uncached ? dirty_3_1 : _GEN_912; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1117 = io_cpu_tlb_uncached ? dirty_4_0 : _GEN_913; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1118 = io_cpu_tlb_uncached ? dirty_4_1 : _GEN_914; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1119 = io_cpu_tlb_uncached ? dirty_5_0 : _GEN_915; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1120 = io_cpu_tlb_uncached ? dirty_5_1 : _GEN_916; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1121 = io_cpu_tlb_uncached ? dirty_6_0 : _GEN_917; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1122 = io_cpu_tlb_uncached ? dirty_6_1 : _GEN_918; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1123 = io_cpu_tlb_uncached ? dirty_7_0 : _GEN_919; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1124 = io_cpu_tlb_uncached ? dirty_7_1 : _GEN_920; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1125 = io_cpu_tlb_uncached ? dirty_8_0 : _GEN_921; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1126 = io_cpu_tlb_uncached ? dirty_8_1 : _GEN_922; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1127 = io_cpu_tlb_uncached ? dirty_9_0 : _GEN_923; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1128 = io_cpu_tlb_uncached ? dirty_9_1 : _GEN_924; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1129 = io_cpu_tlb_uncached ? dirty_10_0 : _GEN_925; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1130 = io_cpu_tlb_uncached ? dirty_10_1 : _GEN_926; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1131 = io_cpu_tlb_uncached ? dirty_11_0 : _GEN_927; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1132 = io_cpu_tlb_uncached ? dirty_11_1 : _GEN_928; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1133 = io_cpu_tlb_uncached ? dirty_12_0 : _GEN_929; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1134 = io_cpu_tlb_uncached ? dirty_12_1 : _GEN_930; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1135 = io_cpu_tlb_uncached ? dirty_13_0 : _GEN_931; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1136 = io_cpu_tlb_uncached ? dirty_13_1 : _GEN_932; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1137 = io_cpu_tlb_uncached ? dirty_14_0 : _GEN_933; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1138 = io_cpu_tlb_uncached ? dirty_14_1 : _GEN_934; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1139 = io_cpu_tlb_uncached ? dirty_15_0 : _GEN_935; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1140 = io_cpu_tlb_uncached ? dirty_15_1 : _GEN_936; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1141 = io_cpu_tlb_uncached ? dirty_16_0 : _GEN_937; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1142 = io_cpu_tlb_uncached ? dirty_16_1 : _GEN_938; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1143 = io_cpu_tlb_uncached ? dirty_17_0 : _GEN_939; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1144 = io_cpu_tlb_uncached ? dirty_17_1 : _GEN_940; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1145 = io_cpu_tlb_uncached ? dirty_18_0 : _GEN_941; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1146 = io_cpu_tlb_uncached ? dirty_18_1 : _GEN_942; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1147 = io_cpu_tlb_uncached ? dirty_19_0 : _GEN_943; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1148 = io_cpu_tlb_uncached ? dirty_19_1 : _GEN_944; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1149 = io_cpu_tlb_uncached ? dirty_20_0 : _GEN_945; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1150 = io_cpu_tlb_uncached ? dirty_20_1 : _GEN_946; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1151 = io_cpu_tlb_uncached ? dirty_21_0 : _GEN_947; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1152 = io_cpu_tlb_uncached ? dirty_21_1 : _GEN_948; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1153 = io_cpu_tlb_uncached ? dirty_22_0 : _GEN_949; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1154 = io_cpu_tlb_uncached ? dirty_22_1 : _GEN_950; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1155 = io_cpu_tlb_uncached ? dirty_23_0 : _GEN_951; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1156 = io_cpu_tlb_uncached ? dirty_23_1 : _GEN_952; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1157 = io_cpu_tlb_uncached ? dirty_24_0 : _GEN_953; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1158 = io_cpu_tlb_uncached ? dirty_24_1 : _GEN_954; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1159 = io_cpu_tlb_uncached ? dirty_25_0 : _GEN_955; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1160 = io_cpu_tlb_uncached ? dirty_25_1 : _GEN_956; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1161 = io_cpu_tlb_uncached ? dirty_26_0 : _GEN_957; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1162 = io_cpu_tlb_uncached ? dirty_26_1 : _GEN_958; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1163 = io_cpu_tlb_uncached ? dirty_27_0 : _GEN_959; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1164 = io_cpu_tlb_uncached ? dirty_27_1 : _GEN_960; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1165 = io_cpu_tlb_uncached ? dirty_28_0 : _GEN_961; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1166 = io_cpu_tlb_uncached ? dirty_28_1 : _GEN_962; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1167 = io_cpu_tlb_uncached ? dirty_29_0 : _GEN_963; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1168 = io_cpu_tlb_uncached ? dirty_29_1 : _GEN_964; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1169 = io_cpu_tlb_uncached ? dirty_30_0 : _GEN_965; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1170 = io_cpu_tlb_uncached ? dirty_30_1 : _GEN_966; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1171 = io_cpu_tlb_uncached ? dirty_31_0 : _GEN_967; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1172 = io_cpu_tlb_uncached ? dirty_31_1 : _GEN_968; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1173 = io_cpu_tlb_uncached ? dirty_32_0 : _GEN_969; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1174 = io_cpu_tlb_uncached ? dirty_32_1 : _GEN_970; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1175 = io_cpu_tlb_uncached ? dirty_33_0 : _GEN_971; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1176 = io_cpu_tlb_uncached ? dirty_33_1 : _GEN_972; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1177 = io_cpu_tlb_uncached ? dirty_34_0 : _GEN_973; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1178 = io_cpu_tlb_uncached ? dirty_34_1 : _GEN_974; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1179 = io_cpu_tlb_uncached ? dirty_35_0 : _GEN_975; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1180 = io_cpu_tlb_uncached ? dirty_35_1 : _GEN_976; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1181 = io_cpu_tlb_uncached ? dirty_36_0 : _GEN_977; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1182 = io_cpu_tlb_uncached ? dirty_36_1 : _GEN_978; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1183 = io_cpu_tlb_uncached ? dirty_37_0 : _GEN_979; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1184 = io_cpu_tlb_uncached ? dirty_37_1 : _GEN_980; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1185 = io_cpu_tlb_uncached ? dirty_38_0 : _GEN_981; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1186 = io_cpu_tlb_uncached ? dirty_38_1 : _GEN_982; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1187 = io_cpu_tlb_uncached ? dirty_39_0 : _GEN_983; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1188 = io_cpu_tlb_uncached ? dirty_39_1 : _GEN_984; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1189 = io_cpu_tlb_uncached ? dirty_40_0 : _GEN_985; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1190 = io_cpu_tlb_uncached ? dirty_40_1 : _GEN_986; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1191 = io_cpu_tlb_uncached ? dirty_41_0 : _GEN_987; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1192 = io_cpu_tlb_uncached ? dirty_41_1 : _GEN_988; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1193 = io_cpu_tlb_uncached ? dirty_42_0 : _GEN_989; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1194 = io_cpu_tlb_uncached ? dirty_42_1 : _GEN_990; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1195 = io_cpu_tlb_uncached ? dirty_43_0 : _GEN_991; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1196 = io_cpu_tlb_uncached ? dirty_43_1 : _GEN_992; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1197 = io_cpu_tlb_uncached ? dirty_44_0 : _GEN_993; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1198 = io_cpu_tlb_uncached ? dirty_44_1 : _GEN_994; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1199 = io_cpu_tlb_uncached ? dirty_45_0 : _GEN_995; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1200 = io_cpu_tlb_uncached ? dirty_45_1 : _GEN_996; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1201 = io_cpu_tlb_uncached ? dirty_46_0 : _GEN_997; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1202 = io_cpu_tlb_uncached ? dirty_46_1 : _GEN_998; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1203 = io_cpu_tlb_uncached ? dirty_47_0 : _GEN_999; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1204 = io_cpu_tlb_uncached ? dirty_47_1 : _GEN_1000; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1205 = io_cpu_tlb_uncached ? dirty_48_0 : _GEN_1001; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1206 = io_cpu_tlb_uncached ? dirty_48_1 : _GEN_1002; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1207 = io_cpu_tlb_uncached ? dirty_49_0 : _GEN_1003; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1208 = io_cpu_tlb_uncached ? dirty_49_1 : _GEN_1004; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1209 = io_cpu_tlb_uncached ? dirty_50_0 : _GEN_1005; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1210 = io_cpu_tlb_uncached ? dirty_50_1 : _GEN_1006; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1211 = io_cpu_tlb_uncached ? dirty_51_0 : _GEN_1007; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1212 = io_cpu_tlb_uncached ? dirty_51_1 : _GEN_1008; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1213 = io_cpu_tlb_uncached ? dirty_52_0 : _GEN_1009; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1214 = io_cpu_tlb_uncached ? dirty_52_1 : _GEN_1010; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1215 = io_cpu_tlb_uncached ? dirty_53_0 : _GEN_1011; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1216 = io_cpu_tlb_uncached ? dirty_53_1 : _GEN_1012; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1217 = io_cpu_tlb_uncached ? dirty_54_0 : _GEN_1013; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1218 = io_cpu_tlb_uncached ? dirty_54_1 : _GEN_1014; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1219 = io_cpu_tlb_uncached ? dirty_55_0 : _GEN_1015; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1220 = io_cpu_tlb_uncached ? dirty_55_1 : _GEN_1016; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1221 = io_cpu_tlb_uncached ? dirty_56_0 : _GEN_1017; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1222 = io_cpu_tlb_uncached ? dirty_56_1 : _GEN_1018; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1223 = io_cpu_tlb_uncached ? dirty_57_0 : _GEN_1019; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1224 = io_cpu_tlb_uncached ? dirty_57_1 : _GEN_1020; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1225 = io_cpu_tlb_uncached ? dirty_58_0 : _GEN_1021; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1226 = io_cpu_tlb_uncached ? dirty_58_1 : _GEN_1022; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1227 = io_cpu_tlb_uncached ? dirty_59_0 : _GEN_1023; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1228 = io_cpu_tlb_uncached ? dirty_59_1 : _GEN_1024; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1229 = io_cpu_tlb_uncached ? dirty_60_0 : _GEN_1025; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1230 = io_cpu_tlb_uncached ? dirty_60_1 : _GEN_1026; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1231 = io_cpu_tlb_uncached ? dirty_61_0 : _GEN_1027; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1232 = io_cpu_tlb_uncached ? dirty_61_1 : _GEN_1028; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1233 = io_cpu_tlb_uncached ? dirty_62_0 : _GEN_1029; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1234 = io_cpu_tlb_uncached ? dirty_62_1 : _GEN_1030; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1235 = io_cpu_tlb_uncached ? dirty_63_0 : _GEN_1031; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire  _GEN_1236 = io_cpu_tlb_uncached ? dirty_63_1 : _GEN_1032; // @[playground/src/cache/DCache.scala 135:22 325:41]
  wire [63:0] _GEN_1237 = io_cpu_tlb_uncached ? saved_rdata : _GEN_1033; // @[playground/src/cache/DCache.scala 209:28 325:41]
  wire [2:0] _GEN_1238 = _dcache_stall_T_3 ? 3'h5 : _GEN_1039; // @[playground/src/cache/DCache.scala 323:37 324:17]
  wire  _GEN_1239 = _dcache_stall_T_3 ? 1'h0 : _GEN_1034; // @[playground/src/cache/DCache.scala 155:26 323:37]
  wire [63:0] _GEN_1240 = _dcache_stall_T_3 ? 64'h0 : _GEN_1035; // @[playground/src/cache/DCache.scala 156:26 323:37]
  wire [7:0] _GEN_1241 = _dcache_stall_T_3 ? 8'h0 : _GEN_1036; // @[playground/src/cache/DCache.scala 156:26 323:37]
  wire [7:0] _GEN_1242 = _dcache_stall_T_3 ? 8'h0 : _GEN_1037; // @[playground/src/cache/DCache.scala 156:26 323:37]
  wire [63:0] _GEN_1243 = _dcache_stall_T_3 ? 64'h0 : _GEN_1038; // @[playground/src/cache/DCache.scala 156:26 323:37]
  wire [31:0] _GEN_1244 = _dcache_stall_T_3 ? ar_addr : _GEN_1040; // @[playground/src/cache/DCache.scala 259:24 323:37]
  wire [7:0] _GEN_1245 = _dcache_stall_T_3 ? ar_len : _GEN_1041; // @[playground/src/cache/DCache.scala 259:24 323:37]
  wire [7:0] _GEN_1246 = _dcache_stall_T_3 ? {{5'd0}, ar_size} : _GEN_1042; // @[playground/src/cache/DCache.scala 259:24 323:37]
  wire  _GEN_1247 = _dcache_stall_T_3 ? arvalid : _GEN_1043; // @[playground/src/cache/DCache.scala 260:24 323:37]
  wire  _GEN_1248 = _dcache_stall_T_3 ? rready : _GEN_1044; // @[playground/src/cache/DCache.scala 263:23 323:37]
  wire  _GEN_1249 = _dcache_stall_T_3 ? lru_0 : _GEN_1045; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1250 = _dcache_stall_T_3 ? lru_1 : _GEN_1046; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1251 = _dcache_stall_T_3 ? lru_2 : _GEN_1047; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1252 = _dcache_stall_T_3 ? lru_3 : _GEN_1048; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1253 = _dcache_stall_T_3 ? lru_4 : _GEN_1049; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1254 = _dcache_stall_T_3 ? lru_5 : _GEN_1050; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1255 = _dcache_stall_T_3 ? lru_6 : _GEN_1051; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1256 = _dcache_stall_T_3 ? lru_7 : _GEN_1052; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1257 = _dcache_stall_T_3 ? lru_8 : _GEN_1053; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1258 = _dcache_stall_T_3 ? lru_9 : _GEN_1054; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1259 = _dcache_stall_T_3 ? lru_10 : _GEN_1055; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1260 = _dcache_stall_T_3 ? lru_11 : _GEN_1056; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1261 = _dcache_stall_T_3 ? lru_12 : _GEN_1057; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1262 = _dcache_stall_T_3 ? lru_13 : _GEN_1058; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1263 = _dcache_stall_T_3 ? lru_14 : _GEN_1059; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1264 = _dcache_stall_T_3 ? lru_15 : _GEN_1060; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1265 = _dcache_stall_T_3 ? lru_16 : _GEN_1061; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1266 = _dcache_stall_T_3 ? lru_17 : _GEN_1062; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1267 = _dcache_stall_T_3 ? lru_18 : _GEN_1063; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1268 = _dcache_stall_T_3 ? lru_19 : _GEN_1064; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1269 = _dcache_stall_T_3 ? lru_20 : _GEN_1065; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1270 = _dcache_stall_T_3 ? lru_21 : _GEN_1066; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1271 = _dcache_stall_T_3 ? lru_22 : _GEN_1067; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1272 = _dcache_stall_T_3 ? lru_23 : _GEN_1068; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1273 = _dcache_stall_T_3 ? lru_24 : _GEN_1069; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1274 = _dcache_stall_T_3 ? lru_25 : _GEN_1070; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1275 = _dcache_stall_T_3 ? lru_26 : _GEN_1071; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1276 = _dcache_stall_T_3 ? lru_27 : _GEN_1072; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1277 = _dcache_stall_T_3 ? lru_28 : _GEN_1073; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1278 = _dcache_stall_T_3 ? lru_29 : _GEN_1074; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1279 = _dcache_stall_T_3 ? lru_30 : _GEN_1075; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1280 = _dcache_stall_T_3 ? lru_31 : _GEN_1076; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1281 = _dcache_stall_T_3 ? lru_32 : _GEN_1077; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1282 = _dcache_stall_T_3 ? lru_33 : _GEN_1078; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1283 = _dcache_stall_T_3 ? lru_34 : _GEN_1079; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1284 = _dcache_stall_T_3 ? lru_35 : _GEN_1080; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1285 = _dcache_stall_T_3 ? lru_36 : _GEN_1081; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1286 = _dcache_stall_T_3 ? lru_37 : _GEN_1082; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1287 = _dcache_stall_T_3 ? lru_38 : _GEN_1083; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1288 = _dcache_stall_T_3 ? lru_39 : _GEN_1084; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1289 = _dcache_stall_T_3 ? lru_40 : _GEN_1085; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1290 = _dcache_stall_T_3 ? lru_41 : _GEN_1086; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1291 = _dcache_stall_T_3 ? lru_42 : _GEN_1087; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1292 = _dcache_stall_T_3 ? lru_43 : _GEN_1088; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1293 = _dcache_stall_T_3 ? lru_44 : _GEN_1089; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1294 = _dcache_stall_T_3 ? lru_45 : _GEN_1090; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1295 = _dcache_stall_T_3 ? lru_46 : _GEN_1091; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1296 = _dcache_stall_T_3 ? lru_47 : _GEN_1092; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1297 = _dcache_stall_T_3 ? lru_48 : _GEN_1093; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1298 = _dcache_stall_T_3 ? lru_49 : _GEN_1094; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1299 = _dcache_stall_T_3 ? lru_50 : _GEN_1095; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1300 = _dcache_stall_T_3 ? lru_51 : _GEN_1096; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1301 = _dcache_stall_T_3 ? lru_52 : _GEN_1097; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1302 = _dcache_stall_T_3 ? lru_53 : _GEN_1098; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1303 = _dcache_stall_T_3 ? lru_54 : _GEN_1099; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1304 = _dcache_stall_T_3 ? lru_55 : _GEN_1100; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1305 = _dcache_stall_T_3 ? lru_56 : _GEN_1101; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1306 = _dcache_stall_T_3 ? lru_57 : _GEN_1102; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1307 = _dcache_stall_T_3 ? lru_58 : _GEN_1103; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1308 = _dcache_stall_T_3 ? lru_59 : _GEN_1104; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1309 = _dcache_stall_T_3 ? lru_60 : _GEN_1105; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1310 = _dcache_stall_T_3 ? lru_61 : _GEN_1106; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1311 = _dcache_stall_T_3 ? lru_62 : _GEN_1107; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1312 = _dcache_stall_T_3 ? lru_63 : _GEN_1108; // @[playground/src/cache/DCache.scala 136:22 323:37]
  wire  _GEN_1313 = _dcache_stall_T_3 ? dirty_0_0 : _GEN_1109; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1314 = _dcache_stall_T_3 ? dirty_0_1 : _GEN_1110; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1315 = _dcache_stall_T_3 ? dirty_1_0 : _GEN_1111; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1316 = _dcache_stall_T_3 ? dirty_1_1 : _GEN_1112; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1317 = _dcache_stall_T_3 ? dirty_2_0 : _GEN_1113; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1318 = _dcache_stall_T_3 ? dirty_2_1 : _GEN_1114; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1319 = _dcache_stall_T_3 ? dirty_3_0 : _GEN_1115; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1320 = _dcache_stall_T_3 ? dirty_3_1 : _GEN_1116; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1321 = _dcache_stall_T_3 ? dirty_4_0 : _GEN_1117; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1322 = _dcache_stall_T_3 ? dirty_4_1 : _GEN_1118; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1323 = _dcache_stall_T_3 ? dirty_5_0 : _GEN_1119; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1324 = _dcache_stall_T_3 ? dirty_5_1 : _GEN_1120; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1325 = _dcache_stall_T_3 ? dirty_6_0 : _GEN_1121; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1326 = _dcache_stall_T_3 ? dirty_6_1 : _GEN_1122; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1327 = _dcache_stall_T_3 ? dirty_7_0 : _GEN_1123; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1328 = _dcache_stall_T_3 ? dirty_7_1 : _GEN_1124; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1329 = _dcache_stall_T_3 ? dirty_8_0 : _GEN_1125; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1330 = _dcache_stall_T_3 ? dirty_8_1 : _GEN_1126; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1331 = _dcache_stall_T_3 ? dirty_9_0 : _GEN_1127; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1332 = _dcache_stall_T_3 ? dirty_9_1 : _GEN_1128; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1333 = _dcache_stall_T_3 ? dirty_10_0 : _GEN_1129; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1334 = _dcache_stall_T_3 ? dirty_10_1 : _GEN_1130; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1335 = _dcache_stall_T_3 ? dirty_11_0 : _GEN_1131; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1336 = _dcache_stall_T_3 ? dirty_11_1 : _GEN_1132; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1337 = _dcache_stall_T_3 ? dirty_12_0 : _GEN_1133; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1338 = _dcache_stall_T_3 ? dirty_12_1 : _GEN_1134; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1339 = _dcache_stall_T_3 ? dirty_13_0 : _GEN_1135; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1340 = _dcache_stall_T_3 ? dirty_13_1 : _GEN_1136; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1341 = _dcache_stall_T_3 ? dirty_14_0 : _GEN_1137; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1342 = _dcache_stall_T_3 ? dirty_14_1 : _GEN_1138; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1343 = _dcache_stall_T_3 ? dirty_15_0 : _GEN_1139; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1344 = _dcache_stall_T_3 ? dirty_15_1 : _GEN_1140; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1345 = _dcache_stall_T_3 ? dirty_16_0 : _GEN_1141; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1346 = _dcache_stall_T_3 ? dirty_16_1 : _GEN_1142; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1347 = _dcache_stall_T_3 ? dirty_17_0 : _GEN_1143; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1348 = _dcache_stall_T_3 ? dirty_17_1 : _GEN_1144; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1349 = _dcache_stall_T_3 ? dirty_18_0 : _GEN_1145; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1350 = _dcache_stall_T_3 ? dirty_18_1 : _GEN_1146; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1351 = _dcache_stall_T_3 ? dirty_19_0 : _GEN_1147; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1352 = _dcache_stall_T_3 ? dirty_19_1 : _GEN_1148; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1353 = _dcache_stall_T_3 ? dirty_20_0 : _GEN_1149; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1354 = _dcache_stall_T_3 ? dirty_20_1 : _GEN_1150; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1355 = _dcache_stall_T_3 ? dirty_21_0 : _GEN_1151; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1356 = _dcache_stall_T_3 ? dirty_21_1 : _GEN_1152; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1357 = _dcache_stall_T_3 ? dirty_22_0 : _GEN_1153; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1358 = _dcache_stall_T_3 ? dirty_22_1 : _GEN_1154; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1359 = _dcache_stall_T_3 ? dirty_23_0 : _GEN_1155; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1360 = _dcache_stall_T_3 ? dirty_23_1 : _GEN_1156; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1361 = _dcache_stall_T_3 ? dirty_24_0 : _GEN_1157; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1362 = _dcache_stall_T_3 ? dirty_24_1 : _GEN_1158; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1363 = _dcache_stall_T_3 ? dirty_25_0 : _GEN_1159; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1364 = _dcache_stall_T_3 ? dirty_25_1 : _GEN_1160; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1365 = _dcache_stall_T_3 ? dirty_26_0 : _GEN_1161; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1366 = _dcache_stall_T_3 ? dirty_26_1 : _GEN_1162; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1367 = _dcache_stall_T_3 ? dirty_27_0 : _GEN_1163; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1368 = _dcache_stall_T_3 ? dirty_27_1 : _GEN_1164; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1369 = _dcache_stall_T_3 ? dirty_28_0 : _GEN_1165; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1370 = _dcache_stall_T_3 ? dirty_28_1 : _GEN_1166; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1371 = _dcache_stall_T_3 ? dirty_29_0 : _GEN_1167; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1372 = _dcache_stall_T_3 ? dirty_29_1 : _GEN_1168; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1373 = _dcache_stall_T_3 ? dirty_30_0 : _GEN_1169; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1374 = _dcache_stall_T_3 ? dirty_30_1 : _GEN_1170; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1375 = _dcache_stall_T_3 ? dirty_31_0 : _GEN_1171; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1376 = _dcache_stall_T_3 ? dirty_31_1 : _GEN_1172; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1377 = _dcache_stall_T_3 ? dirty_32_0 : _GEN_1173; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1378 = _dcache_stall_T_3 ? dirty_32_1 : _GEN_1174; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1379 = _dcache_stall_T_3 ? dirty_33_0 : _GEN_1175; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1380 = _dcache_stall_T_3 ? dirty_33_1 : _GEN_1176; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1381 = _dcache_stall_T_3 ? dirty_34_0 : _GEN_1177; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1382 = _dcache_stall_T_3 ? dirty_34_1 : _GEN_1178; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1383 = _dcache_stall_T_3 ? dirty_35_0 : _GEN_1179; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1384 = _dcache_stall_T_3 ? dirty_35_1 : _GEN_1180; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1385 = _dcache_stall_T_3 ? dirty_36_0 : _GEN_1181; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1386 = _dcache_stall_T_3 ? dirty_36_1 : _GEN_1182; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1387 = _dcache_stall_T_3 ? dirty_37_0 : _GEN_1183; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1388 = _dcache_stall_T_3 ? dirty_37_1 : _GEN_1184; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1389 = _dcache_stall_T_3 ? dirty_38_0 : _GEN_1185; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1390 = _dcache_stall_T_3 ? dirty_38_1 : _GEN_1186; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1391 = _dcache_stall_T_3 ? dirty_39_0 : _GEN_1187; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1392 = _dcache_stall_T_3 ? dirty_39_1 : _GEN_1188; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1393 = _dcache_stall_T_3 ? dirty_40_0 : _GEN_1189; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1394 = _dcache_stall_T_3 ? dirty_40_1 : _GEN_1190; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1395 = _dcache_stall_T_3 ? dirty_41_0 : _GEN_1191; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1396 = _dcache_stall_T_3 ? dirty_41_1 : _GEN_1192; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1397 = _dcache_stall_T_3 ? dirty_42_0 : _GEN_1193; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1398 = _dcache_stall_T_3 ? dirty_42_1 : _GEN_1194; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1399 = _dcache_stall_T_3 ? dirty_43_0 : _GEN_1195; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1400 = _dcache_stall_T_3 ? dirty_43_1 : _GEN_1196; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1401 = _dcache_stall_T_3 ? dirty_44_0 : _GEN_1197; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1402 = _dcache_stall_T_3 ? dirty_44_1 : _GEN_1198; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1403 = _dcache_stall_T_3 ? dirty_45_0 : _GEN_1199; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1404 = _dcache_stall_T_3 ? dirty_45_1 : _GEN_1200; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1405 = _dcache_stall_T_3 ? dirty_46_0 : _GEN_1201; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1406 = _dcache_stall_T_3 ? dirty_46_1 : _GEN_1202; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1407 = _dcache_stall_T_3 ? dirty_47_0 : _GEN_1203; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1408 = _dcache_stall_T_3 ? dirty_47_1 : _GEN_1204; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1409 = _dcache_stall_T_3 ? dirty_48_0 : _GEN_1205; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1410 = _dcache_stall_T_3 ? dirty_48_1 : _GEN_1206; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1411 = _dcache_stall_T_3 ? dirty_49_0 : _GEN_1207; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1412 = _dcache_stall_T_3 ? dirty_49_1 : _GEN_1208; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1413 = _dcache_stall_T_3 ? dirty_50_0 : _GEN_1209; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1414 = _dcache_stall_T_3 ? dirty_50_1 : _GEN_1210; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1415 = _dcache_stall_T_3 ? dirty_51_0 : _GEN_1211; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1416 = _dcache_stall_T_3 ? dirty_51_1 : _GEN_1212; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1417 = _dcache_stall_T_3 ? dirty_52_0 : _GEN_1213; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1418 = _dcache_stall_T_3 ? dirty_52_1 : _GEN_1214; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1419 = _dcache_stall_T_3 ? dirty_53_0 : _GEN_1215; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1420 = _dcache_stall_T_3 ? dirty_53_1 : _GEN_1216; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1421 = _dcache_stall_T_3 ? dirty_54_0 : _GEN_1217; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1422 = _dcache_stall_T_3 ? dirty_54_1 : _GEN_1218; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1423 = _dcache_stall_T_3 ? dirty_55_0 : _GEN_1219; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1424 = _dcache_stall_T_3 ? dirty_55_1 : _GEN_1220; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1425 = _dcache_stall_T_3 ? dirty_56_0 : _GEN_1221; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1426 = _dcache_stall_T_3 ? dirty_56_1 : _GEN_1222; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1427 = _dcache_stall_T_3 ? dirty_57_0 : _GEN_1223; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1428 = _dcache_stall_T_3 ? dirty_57_1 : _GEN_1224; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1429 = _dcache_stall_T_3 ? dirty_58_0 : _GEN_1225; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1430 = _dcache_stall_T_3 ? dirty_58_1 : _GEN_1226; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1431 = _dcache_stall_T_3 ? dirty_59_0 : _GEN_1227; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1432 = _dcache_stall_T_3 ? dirty_59_1 : _GEN_1228; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1433 = _dcache_stall_T_3 ? dirty_60_0 : _GEN_1229; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1434 = _dcache_stall_T_3 ? dirty_60_1 : _GEN_1230; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1435 = _dcache_stall_T_3 ? dirty_61_0 : _GEN_1231; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1436 = _dcache_stall_T_3 ? dirty_61_1 : _GEN_1232; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1437 = _dcache_stall_T_3 ? dirty_62_0 : _GEN_1233; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1438 = _dcache_stall_T_3 ? dirty_62_1 : _GEN_1234; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1439 = _dcache_stall_T_3 ? dirty_63_0 : _GEN_1235; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire  _GEN_1440 = _dcache_stall_T_3 ? dirty_63_1 : _GEN_1236; // @[playground/src/cache/DCache.scala 135:22 323:37]
  wire [63:0] _GEN_1441 = _dcache_stall_T_3 ? saved_rdata : _GEN_1237; // @[playground/src/cache/DCache.scala 209:28 323:37]
  wire [2:0] _GEN_1443 = addr_err ? state : _GEN_1238; // @[playground/src/cache/DCache.scala 321:24 90:94]
  wire  _GEN_1444 = addr_err ? 1'h0 : _GEN_1239; // @[playground/src/cache/DCache.scala 321:24 155:26]
  wire [63:0] _GEN_1445 = addr_err ? 64'h0 : _GEN_1240; // @[playground/src/cache/DCache.scala 321:24 156:26]
  wire [7:0] _GEN_1446 = addr_err ? 8'h0 : _GEN_1241; // @[playground/src/cache/DCache.scala 321:24 156:26]
  wire [7:0] _GEN_1447 = addr_err ? 8'h0 : _GEN_1242; // @[playground/src/cache/DCache.scala 321:24 156:26]
  wire [63:0] _GEN_1448 = addr_err ? 64'h0 : _GEN_1243; // @[playground/src/cache/DCache.scala 321:24 156:26]
  wire [31:0] _GEN_1449 = addr_err ? ar_addr : _GEN_1244; // @[playground/src/cache/DCache.scala 259:24 321:24]
  wire [7:0] _GEN_1450 = addr_err ? ar_len : _GEN_1245; // @[playground/src/cache/DCache.scala 259:24 321:24]
  wire [7:0] _GEN_1451 = addr_err ? {{5'd0}, ar_size} : _GEN_1246; // @[playground/src/cache/DCache.scala 259:24 321:24]
  wire  _GEN_1452 = addr_err ? arvalid : _GEN_1247; // @[playground/src/cache/DCache.scala 260:24 321:24]
  wire  _GEN_1453 = addr_err ? rready : _GEN_1248; // @[playground/src/cache/DCache.scala 263:23 321:24]
  wire  _io_cpu_tlb_ptw_vpn_ready_T = ~ptw_working; // @[playground/src/cache/DCache.scala 364:37]
  wire [7:0] lo_lo_lo_lo = {dirty_3_1,dirty_3_0,dirty_2_1,dirty_2_0,dirty_1_1,dirty_1_0,dirty_0_1,dirty_0_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [15:0] lo_lo_lo = {dirty_7_1,dirty_7_0,dirty_6_1,dirty_6_0,dirty_5_1,dirty_5_0,dirty_4_1,dirty_4_0,lo_lo_lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] lo_lo_hi_lo = {dirty_11_1,dirty_11_0,dirty_10_1,dirty_10_0,dirty_9_1,dirty_9_0,dirty_8_1,dirty_8_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [31:0] lo_lo = {dirty_15_1,dirty_15_0,dirty_14_1,dirty_14_0,dirty_13_1,dirty_13_0,dirty_12_1,dirty_12_0,
    lo_lo_hi_lo,lo_lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] lo_hi_lo_lo = {dirty_19_1,dirty_19_0,dirty_18_1,dirty_18_0,dirty_17_1,dirty_17_0,dirty_16_1,dirty_16_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [15:0] lo_hi_lo = {dirty_23_1,dirty_23_0,dirty_22_1,dirty_22_0,dirty_21_1,dirty_21_0,dirty_20_1,dirty_20_0,
    lo_hi_lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] lo_hi_hi_lo = {dirty_27_1,dirty_27_0,dirty_26_1,dirty_26_0,dirty_25_1,dirty_25_0,dirty_24_1,dirty_24_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [31:0] lo_hi = {dirty_31_1,dirty_31_0,dirty_30_1,dirty_30_0,dirty_29_1,dirty_29_0,dirty_28_1,dirty_28_0,
    lo_hi_hi_lo,lo_hi_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] hi_lo_lo_lo = {dirty_35_1,dirty_35_0,dirty_34_1,dirty_34_0,dirty_33_1,dirty_33_0,dirty_32_1,dirty_32_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [15:0] hi_lo_lo = {dirty_39_1,dirty_39_0,dirty_38_1,dirty_38_0,dirty_37_1,dirty_37_0,dirty_36_1,dirty_36_0,
    hi_lo_lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] hi_lo_hi_lo = {dirty_43_1,dirty_43_0,dirty_42_1,dirty_42_0,dirty_41_1,dirty_41_0,dirty_40_1,dirty_40_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [31:0] hi_lo = {dirty_47_1,dirty_47_0,dirty_46_1,dirty_46_0,dirty_45_1,dirty_45_0,dirty_44_1,dirty_44_0,
    hi_lo_hi_lo,hi_lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] hi_hi_lo_lo = {dirty_51_1,dirty_51_0,dirty_50_1,dirty_50_0,dirty_49_1,dirty_49_0,dirty_48_1,dirty_48_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [15:0] hi_hi_lo = {dirty_55_1,dirty_55_0,dirty_54_1,dirty_54_0,dirty_53_1,dirty_53_0,dirty_52_1,dirty_52_0,
    hi_hi_lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [7:0] hi_hi_hi_lo = {dirty_59_1,dirty_59_0,dirty_58_1,dirty_58_0,dirty_57_1,dirty_57_0,dirty_56_1,dirty_56_0}; // @[playground/src/cache/DCache.scala 367:22]
  wire [31:0] hi_hi = {dirty_63_1,dirty_63_0,dirty_62_1,dirty_62_0,dirty_61_1,dirty_61_0,dirty_60_1,dirty_60_0,
    hi_hi_hi_lo,hi_hi_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire [127:0] _T_13 = {hi_hi,hi_lo,lo_hi,lo_lo}; // @[playground/src/cache/DCache.scala 367:22]
  wire  _T_14 = |_T_13; // @[playground/src/cache/DCache.scala 367:29]
  wire [2:0] _GEN_1647 = _T_8 ? 3'h2 : state; // @[playground/src/cache/DCache.scala 368:35 369:24 90:94]
  wire  _GEN_1648 = _T_8 ? 1'h0 : readsram; // @[playground/src/cache/DCache.scala 368:35 370:24 148:25]
  wire [2:0] _GEN_1649 = |_T_13 ? _GEN_1647 : 3'h4; // @[playground/src/cache/DCache.scala 367:34 374:19]
  wire  _GEN_1650 = |_T_13 ? _GEN_1648 : readsram; // @[playground/src/cache/DCache.scala 148:25 367:34]
  wire [2:0] _GEN_1651 = io_cpu_fence_i ? _GEN_1649 : state; // @[playground/src/cache/DCache.scala 365:30 90:94]
  wire  _GEN_1653 = io_cpu_en & addr_err; // @[playground/src/cache/DCache.scala 318:20 320:23]
  wire [2:0] _GEN_1654 = io_cpu_en ? _GEN_1443 : _GEN_1651; // @[playground/src/cache/DCache.scala 320:23]
  wire  _GEN_1655 = io_cpu_en & _GEN_1444; // @[playground/src/cache/DCache.scala 320:23 155:26]
  wire [63:0] _GEN_1656 = io_cpu_en ? _GEN_1445 : 64'h0; // @[playground/src/cache/DCache.scala 320:23 156:26]
  wire [7:0] _GEN_1657 = io_cpu_en ? _GEN_1446 : 8'h0; // @[playground/src/cache/DCache.scala 320:23 156:26]
  wire [7:0] _GEN_1658 = io_cpu_en ? _GEN_1447 : 8'h0; // @[playground/src/cache/DCache.scala 320:23 156:26]
  wire [63:0] _GEN_1659 = io_cpu_en ? _GEN_1448 : 64'h0; // @[playground/src/cache/DCache.scala 320:23 156:26]
  wire [31:0] _GEN_1660 = io_cpu_en ? _GEN_1449 : ar_addr; // @[playground/src/cache/DCache.scala 320:23 259:24]
  wire [7:0] _GEN_1661 = io_cpu_en ? _GEN_1450 : ar_len; // @[playground/src/cache/DCache.scala 320:23 259:24]
  wire [7:0] _GEN_1662 = io_cpu_en ? _GEN_1451 : {{5'd0}, ar_size}; // @[playground/src/cache/DCache.scala 320:23 259:24]
  wire  _GEN_1663 = io_cpu_en ? _GEN_1452 : arvalid; // @[playground/src/cache/DCache.scala 320:23 260:24]
  wire  _GEN_1664 = io_cpu_en ? _GEN_1453 : rready; // @[playground/src/cache/DCache.scala 263:23 320:23]
  wire  _GEN_1858 = io_cpu_en ? 1'h0 : ~ptw_working; // @[playground/src/cache/DCache.scala 320:23 107:28 364:34]
  wire  _GEN_1860 = arvalid & io_axi_ar_ready ? 1'h0 : arvalid; // @[playground/src/cache/DCache.scala 380:40 381:17 260:24]
  wire  _T_18 = io_axi_r_ready & io_axi_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _GEN_1861 = _T_18 ? 1'h0 : rready; // @[playground/src/cache/DCache.scala 383:27 384:22 263:23]
  wire [2:0] _GEN_1864 = _T_18 ? 3'h4 : state; // @[playground/src/cache/DCache.scala 383:27 387:22 90:94]
  wire  _GEN_1865 = _T ? 1'h0 : _GEN_290; // @[playground/src/cache/DCache.scala 392:30 393:19]
  wire [2:0] _bank_wbindex_T_1 = bank_wbindex + 3'h1; // @[playground/src/cache/DCache.scala 399:42]
  wire  _GEN_1867 = 6'h1 == dirty_index ? dirty_1_1 : dirty_0_1; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1868 = 6'h2 == dirty_index ? dirty_2_1 : _GEN_1867; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1869 = 6'h3 == dirty_index ? dirty_3_1 : _GEN_1868; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1870 = 6'h4 == dirty_index ? dirty_4_1 : _GEN_1869; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1871 = 6'h5 == dirty_index ? dirty_5_1 : _GEN_1870; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1872 = 6'h6 == dirty_index ? dirty_6_1 : _GEN_1871; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1873 = 6'h7 == dirty_index ? dirty_7_1 : _GEN_1872; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1874 = 6'h8 == dirty_index ? dirty_8_1 : _GEN_1873; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1875 = 6'h9 == dirty_index ? dirty_9_1 : _GEN_1874; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1876 = 6'ha == dirty_index ? dirty_10_1 : _GEN_1875; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1877 = 6'hb == dirty_index ? dirty_11_1 : _GEN_1876; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1878 = 6'hc == dirty_index ? dirty_12_1 : _GEN_1877; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1879 = 6'hd == dirty_index ? dirty_13_1 : _GEN_1878; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1880 = 6'he == dirty_index ? dirty_14_1 : _GEN_1879; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1881 = 6'hf == dirty_index ? dirty_15_1 : _GEN_1880; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1882 = 6'h10 == dirty_index ? dirty_16_1 : _GEN_1881; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1883 = 6'h11 == dirty_index ? dirty_17_1 : _GEN_1882; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1884 = 6'h12 == dirty_index ? dirty_18_1 : _GEN_1883; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1885 = 6'h13 == dirty_index ? dirty_19_1 : _GEN_1884; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1886 = 6'h14 == dirty_index ? dirty_20_1 : _GEN_1885; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1887 = 6'h15 == dirty_index ? dirty_21_1 : _GEN_1886; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1888 = 6'h16 == dirty_index ? dirty_22_1 : _GEN_1887; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1889 = 6'h17 == dirty_index ? dirty_23_1 : _GEN_1888; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1890 = 6'h18 == dirty_index ? dirty_24_1 : _GEN_1889; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1891 = 6'h19 == dirty_index ? dirty_25_1 : _GEN_1890; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1892 = 6'h1a == dirty_index ? dirty_26_1 : _GEN_1891; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1893 = 6'h1b == dirty_index ? dirty_27_1 : _GEN_1892; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1894 = 6'h1c == dirty_index ? dirty_28_1 : _GEN_1893; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1895 = 6'h1d == dirty_index ? dirty_29_1 : _GEN_1894; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1896 = 6'h1e == dirty_index ? dirty_30_1 : _GEN_1895; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1897 = 6'h1f == dirty_index ? dirty_31_1 : _GEN_1896; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1898 = 6'h20 == dirty_index ? dirty_32_1 : _GEN_1897; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1899 = 6'h21 == dirty_index ? dirty_33_1 : _GEN_1898; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1900 = 6'h22 == dirty_index ? dirty_34_1 : _GEN_1899; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1901 = 6'h23 == dirty_index ? dirty_35_1 : _GEN_1900; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1902 = 6'h24 == dirty_index ? dirty_36_1 : _GEN_1901; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1903 = 6'h25 == dirty_index ? dirty_37_1 : _GEN_1902; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1904 = 6'h26 == dirty_index ? dirty_38_1 : _GEN_1903; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1905 = 6'h27 == dirty_index ? dirty_39_1 : _GEN_1904; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1906 = 6'h28 == dirty_index ? dirty_40_1 : _GEN_1905; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1907 = 6'h29 == dirty_index ? dirty_41_1 : _GEN_1906; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1908 = 6'h2a == dirty_index ? dirty_42_1 : _GEN_1907; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1909 = 6'h2b == dirty_index ? dirty_43_1 : _GEN_1908; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1910 = 6'h2c == dirty_index ? dirty_44_1 : _GEN_1909; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1911 = 6'h2d == dirty_index ? dirty_45_1 : _GEN_1910; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1912 = 6'h2e == dirty_index ? dirty_46_1 : _GEN_1911; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1913 = 6'h2f == dirty_index ? dirty_47_1 : _GEN_1912; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1914 = 6'h30 == dirty_index ? dirty_48_1 : _GEN_1913; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1915 = 6'h31 == dirty_index ? dirty_49_1 : _GEN_1914; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1916 = 6'h32 == dirty_index ? dirty_50_1 : _GEN_1915; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1917 = 6'h33 == dirty_index ? dirty_51_1 : _GEN_1916; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1918 = 6'h34 == dirty_index ? dirty_52_1 : _GEN_1917; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1919 = 6'h35 == dirty_index ? dirty_53_1 : _GEN_1918; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1920 = 6'h36 == dirty_index ? dirty_54_1 : _GEN_1919; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1921 = 6'h37 == dirty_index ? dirty_55_1 : _GEN_1920; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1922 = 6'h38 == dirty_index ? dirty_56_1 : _GEN_1921; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1923 = 6'h39 == dirty_index ? dirty_57_1 : _GEN_1922; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1924 = 6'h3a == dirty_index ? dirty_58_1 : _GEN_1923; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1925 = 6'h3b == dirty_index ? dirty_59_1 : _GEN_1924; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1926 = 6'h3c == dirty_index ? dirty_60_1 : _GEN_1925; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1927 = 6'h3d == dirty_index ? dirty_61_1 : _GEN_1926; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1928 = 6'h3e == dirty_index ? dirty_62_1 : _GEN_1927; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1929 = 6'h3f == dirty_index ? dirty_63_1 : _GEN_1928; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1931 = 3'h0 == _bank_wbindex_T_1 & _GEN_1929 ? data_0_1 : data_0_0; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_6610 = ~_GEN_1929; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1932 = 3'h1 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_1_0 : _GEN_1931; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1933 = 3'h1 == _bank_wbindex_T_1 & _GEN_1929 ? data_1_1 : _GEN_1932; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1934 = 3'h2 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_2_0 : _GEN_1933; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1935 = 3'h2 == _bank_wbindex_T_1 & _GEN_1929 ? data_2_1 : _GEN_1934; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1936 = 3'h3 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_3_0 : _GEN_1935; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1937 = 3'h3 == _bank_wbindex_T_1 & _GEN_1929 ? data_3_1 : _GEN_1936; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1938 = 3'h4 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_4_0 : _GEN_1937; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1939 = 3'h4 == _bank_wbindex_T_1 & _GEN_1929 ? data_4_1 : _GEN_1938; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1940 = 3'h5 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_5_0 : _GEN_1939; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1941 = 3'h5 == _bank_wbindex_T_1 & _GEN_1929 ? data_5_1 : _GEN_1940; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1942 = 3'h6 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_6_0 : _GEN_1941; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1943 = 3'h6 == _bank_wbindex_T_1 & _GEN_1929 ? data_6_1 : _GEN_1942; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1944 = 3'h7 == _bank_wbindex_T_1 & ~_GEN_1929 ? data_7_0 : _GEN_1943; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire [63:0] _GEN_1945 = 3'h7 == _bank_wbindex_T_1 & _GEN_1929 ? data_7_1 : _GEN_1944; // @[playground/src/cache/DCache.scala 400:{26,26}]
  wire  _GEN_1946 = _bank_wbindex_T_1 == 3'h7 | _GEN_292; // @[playground/src/cache/DCache.scala 401:57 402:22]
  wire  _GEN_1947 = w_last ? 1'h0 : _GEN_291; // @[playground/src/cache/DCache.scala 396:24 397:20]
  wire [2:0] _GEN_1948 = w_last ? bank_wbindex : _bank_wbindex_T_1; // @[playground/src/cache/DCache.scala 396:24 165:29 399:26]
  wire [63:0] _GEN_1949 = w_last ? _GEN_297 : _GEN_1945; // @[playground/src/cache/DCache.scala 396:24 400:26]
  wire  _GEN_1950 = w_last ? _GEN_292 : _GEN_1946; // @[playground/src/cache/DCache.scala 396:24]
  wire  _GEN_1951 = _T_1 ? _GEN_1947 : _GEN_291; // @[playground/src/cache/DCache.scala 395:29]
  wire [2:0] _GEN_1952 = _T_1 ? _GEN_1948 : bank_wbindex; // @[playground/src/cache/DCache.scala 165:29 395:29]
  wire [63:0] _GEN_1953 = _T_1 ? _GEN_1949 : _GEN_297; // @[playground/src/cache/DCache.scala 395:29]
  wire  _GEN_1954 = _T_1 ? _GEN_1950 : _GEN_292; // @[playground/src/cache/DCache.scala 395:29]
  wire  _GEN_1955 = 6'h0 == dirty_index & _GEN_6610 ? 1'h0 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1956 = 6'h0 == dirty_index & _GEN_1929 ? 1'h0 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1957 = 6'h1 == dirty_index & _GEN_6610 ? 1'h0 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1958 = 6'h1 == dirty_index & _GEN_1929 ? 1'h0 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1959 = 6'h2 == dirty_index & _GEN_6610 ? 1'h0 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1960 = 6'h2 == dirty_index & _GEN_1929 ? 1'h0 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1961 = 6'h3 == dirty_index & _GEN_6610 ? 1'h0 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1962 = 6'h3 == dirty_index & _GEN_1929 ? 1'h0 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1963 = 6'h4 == dirty_index & _GEN_6610 ? 1'h0 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1964 = 6'h4 == dirty_index & _GEN_1929 ? 1'h0 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1965 = 6'h5 == dirty_index & _GEN_6610 ? 1'h0 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1966 = 6'h5 == dirty_index & _GEN_1929 ? 1'h0 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1967 = 6'h6 == dirty_index & _GEN_6610 ? 1'h0 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1968 = 6'h6 == dirty_index & _GEN_1929 ? 1'h0 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1969 = 6'h7 == dirty_index & _GEN_6610 ? 1'h0 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1970 = 6'h7 == dirty_index & _GEN_1929 ? 1'h0 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1971 = 6'h8 == dirty_index & _GEN_6610 ? 1'h0 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1972 = 6'h8 == dirty_index & _GEN_1929 ? 1'h0 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1973 = 6'h9 == dirty_index & _GEN_6610 ? 1'h0 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1974 = 6'h9 == dirty_index & _GEN_1929 ? 1'h0 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1975 = 6'ha == dirty_index & _GEN_6610 ? 1'h0 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1976 = 6'ha == dirty_index & _GEN_1929 ? 1'h0 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1977 = 6'hb == dirty_index & _GEN_6610 ? 1'h0 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1978 = 6'hb == dirty_index & _GEN_1929 ? 1'h0 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1979 = 6'hc == dirty_index & _GEN_6610 ? 1'h0 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1980 = 6'hc == dirty_index & _GEN_1929 ? 1'h0 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1981 = 6'hd == dirty_index & _GEN_6610 ? 1'h0 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1982 = 6'hd == dirty_index & _GEN_1929 ? 1'h0 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1983 = 6'he == dirty_index & _GEN_6610 ? 1'h0 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1984 = 6'he == dirty_index & _GEN_1929 ? 1'h0 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1985 = 6'hf == dirty_index & _GEN_6610 ? 1'h0 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1986 = 6'hf == dirty_index & _GEN_1929 ? 1'h0 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1987 = 6'h10 == dirty_index & _GEN_6610 ? 1'h0 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1988 = 6'h10 == dirty_index & _GEN_1929 ? 1'h0 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1989 = 6'h11 == dirty_index & _GEN_6610 ? 1'h0 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1990 = 6'h11 == dirty_index & _GEN_1929 ? 1'h0 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1991 = 6'h12 == dirty_index & _GEN_6610 ? 1'h0 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1992 = 6'h12 == dirty_index & _GEN_1929 ? 1'h0 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1993 = 6'h13 == dirty_index & _GEN_6610 ? 1'h0 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1994 = 6'h13 == dirty_index & _GEN_1929 ? 1'h0 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1995 = 6'h14 == dirty_index & _GEN_6610 ? 1'h0 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1996 = 6'h14 == dirty_index & _GEN_1929 ? 1'h0 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1997 = 6'h15 == dirty_index & _GEN_6610 ? 1'h0 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1998 = 6'h15 == dirty_index & _GEN_1929 ? 1'h0 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_1999 = 6'h16 == dirty_index & _GEN_6610 ? 1'h0 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2000 = 6'h16 == dirty_index & _GEN_1929 ? 1'h0 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2001 = 6'h17 == dirty_index & _GEN_6610 ? 1'h0 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2002 = 6'h17 == dirty_index & _GEN_1929 ? 1'h0 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2003 = 6'h18 == dirty_index & _GEN_6610 ? 1'h0 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2004 = 6'h18 == dirty_index & _GEN_1929 ? 1'h0 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2005 = 6'h19 == dirty_index & _GEN_6610 ? 1'h0 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2006 = 6'h19 == dirty_index & _GEN_1929 ? 1'h0 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2007 = 6'h1a == dirty_index & _GEN_6610 ? 1'h0 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2008 = 6'h1a == dirty_index & _GEN_1929 ? 1'h0 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2009 = 6'h1b == dirty_index & _GEN_6610 ? 1'h0 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2010 = 6'h1b == dirty_index & _GEN_1929 ? 1'h0 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2011 = 6'h1c == dirty_index & _GEN_6610 ? 1'h0 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2012 = 6'h1c == dirty_index & _GEN_1929 ? 1'h0 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2013 = 6'h1d == dirty_index & _GEN_6610 ? 1'h0 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2014 = 6'h1d == dirty_index & _GEN_1929 ? 1'h0 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2015 = 6'h1e == dirty_index & _GEN_6610 ? 1'h0 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2016 = 6'h1e == dirty_index & _GEN_1929 ? 1'h0 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2017 = 6'h1f == dirty_index & _GEN_6610 ? 1'h0 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2018 = 6'h1f == dirty_index & _GEN_1929 ? 1'h0 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2019 = 6'h20 == dirty_index & _GEN_6610 ? 1'h0 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2020 = 6'h20 == dirty_index & _GEN_1929 ? 1'h0 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2021 = 6'h21 == dirty_index & _GEN_6610 ? 1'h0 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2022 = 6'h21 == dirty_index & _GEN_1929 ? 1'h0 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2023 = 6'h22 == dirty_index & _GEN_6610 ? 1'h0 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2024 = 6'h22 == dirty_index & _GEN_1929 ? 1'h0 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2025 = 6'h23 == dirty_index & _GEN_6610 ? 1'h0 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2026 = 6'h23 == dirty_index & _GEN_1929 ? 1'h0 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2027 = 6'h24 == dirty_index & _GEN_6610 ? 1'h0 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2028 = 6'h24 == dirty_index & _GEN_1929 ? 1'h0 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2029 = 6'h25 == dirty_index & _GEN_6610 ? 1'h0 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2030 = 6'h25 == dirty_index & _GEN_1929 ? 1'h0 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2031 = 6'h26 == dirty_index & _GEN_6610 ? 1'h0 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2032 = 6'h26 == dirty_index & _GEN_1929 ? 1'h0 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2033 = 6'h27 == dirty_index & _GEN_6610 ? 1'h0 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2034 = 6'h27 == dirty_index & _GEN_1929 ? 1'h0 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2035 = 6'h28 == dirty_index & _GEN_6610 ? 1'h0 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2036 = 6'h28 == dirty_index & _GEN_1929 ? 1'h0 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2037 = 6'h29 == dirty_index & _GEN_6610 ? 1'h0 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2038 = 6'h29 == dirty_index & _GEN_1929 ? 1'h0 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2039 = 6'h2a == dirty_index & _GEN_6610 ? 1'h0 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2040 = 6'h2a == dirty_index & _GEN_1929 ? 1'h0 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2041 = 6'h2b == dirty_index & _GEN_6610 ? 1'h0 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2042 = 6'h2b == dirty_index & _GEN_1929 ? 1'h0 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2043 = 6'h2c == dirty_index & _GEN_6610 ? 1'h0 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2044 = 6'h2c == dirty_index & _GEN_1929 ? 1'h0 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2045 = 6'h2d == dirty_index & _GEN_6610 ? 1'h0 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2046 = 6'h2d == dirty_index & _GEN_1929 ? 1'h0 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2047 = 6'h2e == dirty_index & _GEN_6610 ? 1'h0 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2048 = 6'h2e == dirty_index & _GEN_1929 ? 1'h0 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2049 = 6'h2f == dirty_index & _GEN_6610 ? 1'h0 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2050 = 6'h2f == dirty_index & _GEN_1929 ? 1'h0 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2051 = 6'h30 == dirty_index & _GEN_6610 ? 1'h0 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2052 = 6'h30 == dirty_index & _GEN_1929 ? 1'h0 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2053 = 6'h31 == dirty_index & _GEN_6610 ? 1'h0 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2054 = 6'h31 == dirty_index & _GEN_1929 ? 1'h0 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2055 = 6'h32 == dirty_index & _GEN_6610 ? 1'h0 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2056 = 6'h32 == dirty_index & _GEN_1929 ? 1'h0 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2057 = 6'h33 == dirty_index & _GEN_6610 ? 1'h0 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2058 = 6'h33 == dirty_index & _GEN_1929 ? 1'h0 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2059 = 6'h34 == dirty_index & _GEN_6610 ? 1'h0 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2060 = 6'h34 == dirty_index & _GEN_1929 ? 1'h0 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2061 = 6'h35 == dirty_index & _GEN_6610 ? 1'h0 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2062 = 6'h35 == dirty_index & _GEN_1929 ? 1'h0 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2063 = 6'h36 == dirty_index & _GEN_6610 ? 1'h0 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2064 = 6'h36 == dirty_index & _GEN_1929 ? 1'h0 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2065 = 6'h37 == dirty_index & _GEN_6610 ? 1'h0 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2066 = 6'h37 == dirty_index & _GEN_1929 ? 1'h0 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2067 = 6'h38 == dirty_index & _GEN_6610 ? 1'h0 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2068 = 6'h38 == dirty_index & _GEN_1929 ? 1'h0 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2069 = 6'h39 == dirty_index & _GEN_6610 ? 1'h0 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2070 = 6'h39 == dirty_index & _GEN_1929 ? 1'h0 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2071 = 6'h3a == dirty_index & _GEN_6610 ? 1'h0 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2072 = 6'h3a == dirty_index & _GEN_1929 ? 1'h0 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2073 = 6'h3b == dirty_index & _GEN_6610 ? 1'h0 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2074 = 6'h3b == dirty_index & _GEN_1929 ? 1'h0 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2075 = 6'h3c == dirty_index & _GEN_6610 ? 1'h0 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2076 = 6'h3c == dirty_index & _GEN_1929 ? 1'h0 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2077 = 6'h3d == dirty_index & _GEN_6610 ? 1'h0 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2078 = 6'h3d == dirty_index & _GEN_1929 ? 1'h0 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2079 = 6'h3e == dirty_index & _GEN_6610 ? 1'h0 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2080 = 6'h3e == dirty_index & _GEN_1929 ? 1'h0 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2081 = 6'h3f == dirty_index & _GEN_6610 ? 1'h0 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2082 = 6'h3f == dirty_index & _GEN_1929 ? 1'h0 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 409:{41,41}]
  wire  _GEN_2083 = io_axi_b_valid ? _GEN_1955 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2084 = io_axi_b_valid ? _GEN_1956 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2085 = io_axi_b_valid ? _GEN_1957 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2086 = io_axi_b_valid ? _GEN_1958 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2087 = io_axi_b_valid ? _GEN_1959 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2088 = io_axi_b_valid ? _GEN_1960 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2089 = io_axi_b_valid ? _GEN_1961 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2090 = io_axi_b_valid ? _GEN_1962 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2091 = io_axi_b_valid ? _GEN_1963 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2092 = io_axi_b_valid ? _GEN_1964 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2093 = io_axi_b_valid ? _GEN_1965 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2094 = io_axi_b_valid ? _GEN_1966 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2095 = io_axi_b_valid ? _GEN_1967 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2096 = io_axi_b_valid ? _GEN_1968 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2097 = io_axi_b_valid ? _GEN_1969 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2098 = io_axi_b_valid ? _GEN_1970 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2099 = io_axi_b_valid ? _GEN_1971 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2100 = io_axi_b_valid ? _GEN_1972 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2101 = io_axi_b_valid ? _GEN_1973 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2102 = io_axi_b_valid ? _GEN_1974 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2103 = io_axi_b_valid ? _GEN_1975 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2104 = io_axi_b_valid ? _GEN_1976 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2105 = io_axi_b_valid ? _GEN_1977 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2106 = io_axi_b_valid ? _GEN_1978 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2107 = io_axi_b_valid ? _GEN_1979 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2108 = io_axi_b_valid ? _GEN_1980 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2109 = io_axi_b_valid ? _GEN_1981 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2110 = io_axi_b_valid ? _GEN_1982 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2111 = io_axi_b_valid ? _GEN_1983 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2112 = io_axi_b_valid ? _GEN_1984 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2113 = io_axi_b_valid ? _GEN_1985 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2114 = io_axi_b_valid ? _GEN_1986 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2115 = io_axi_b_valid ? _GEN_1987 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2116 = io_axi_b_valid ? _GEN_1988 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2117 = io_axi_b_valid ? _GEN_1989 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2118 = io_axi_b_valid ? _GEN_1990 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2119 = io_axi_b_valid ? _GEN_1991 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2120 = io_axi_b_valid ? _GEN_1992 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2121 = io_axi_b_valid ? _GEN_1993 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2122 = io_axi_b_valid ? _GEN_1994 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2123 = io_axi_b_valid ? _GEN_1995 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2124 = io_axi_b_valid ? _GEN_1996 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2125 = io_axi_b_valid ? _GEN_1997 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2126 = io_axi_b_valid ? _GEN_1998 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2127 = io_axi_b_valid ? _GEN_1999 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2128 = io_axi_b_valid ? _GEN_2000 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2129 = io_axi_b_valid ? _GEN_2001 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2130 = io_axi_b_valid ? _GEN_2002 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2131 = io_axi_b_valid ? _GEN_2003 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2132 = io_axi_b_valid ? _GEN_2004 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2133 = io_axi_b_valid ? _GEN_2005 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2134 = io_axi_b_valid ? _GEN_2006 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2135 = io_axi_b_valid ? _GEN_2007 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2136 = io_axi_b_valid ? _GEN_2008 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2137 = io_axi_b_valid ? _GEN_2009 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2138 = io_axi_b_valid ? _GEN_2010 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2139 = io_axi_b_valid ? _GEN_2011 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2140 = io_axi_b_valid ? _GEN_2012 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2141 = io_axi_b_valid ? _GEN_2013 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2142 = io_axi_b_valid ? _GEN_2014 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2143 = io_axi_b_valid ? _GEN_2015 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2144 = io_axi_b_valid ? _GEN_2016 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2145 = io_axi_b_valid ? _GEN_2017 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2146 = io_axi_b_valid ? _GEN_2018 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2147 = io_axi_b_valid ? _GEN_2019 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2148 = io_axi_b_valid ? _GEN_2020 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2149 = io_axi_b_valid ? _GEN_2021 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2150 = io_axi_b_valid ? _GEN_2022 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2151 = io_axi_b_valid ? _GEN_2023 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2152 = io_axi_b_valid ? _GEN_2024 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2153 = io_axi_b_valid ? _GEN_2025 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2154 = io_axi_b_valid ? _GEN_2026 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2155 = io_axi_b_valid ? _GEN_2027 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2156 = io_axi_b_valid ? _GEN_2028 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2157 = io_axi_b_valid ? _GEN_2029 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2158 = io_axi_b_valid ? _GEN_2030 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2159 = io_axi_b_valid ? _GEN_2031 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2160 = io_axi_b_valid ? _GEN_2032 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2161 = io_axi_b_valid ? _GEN_2033 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2162 = io_axi_b_valid ? _GEN_2034 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2163 = io_axi_b_valid ? _GEN_2035 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2164 = io_axi_b_valid ? _GEN_2036 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2165 = io_axi_b_valid ? _GEN_2037 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2166 = io_axi_b_valid ? _GEN_2038 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2167 = io_axi_b_valid ? _GEN_2039 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2168 = io_axi_b_valid ? _GEN_2040 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2169 = io_axi_b_valid ? _GEN_2041 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2170 = io_axi_b_valid ? _GEN_2042 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2171 = io_axi_b_valid ? _GEN_2043 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2172 = io_axi_b_valid ? _GEN_2044 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2173 = io_axi_b_valid ? _GEN_2045 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2174 = io_axi_b_valid ? _GEN_2046 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2175 = io_axi_b_valid ? _GEN_2047 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2176 = io_axi_b_valid ? _GEN_2048 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2177 = io_axi_b_valid ? _GEN_2049 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2178 = io_axi_b_valid ? _GEN_2050 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2179 = io_axi_b_valid ? _GEN_2051 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2180 = io_axi_b_valid ? _GEN_2052 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2181 = io_axi_b_valid ? _GEN_2053 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2182 = io_axi_b_valid ? _GEN_2054 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2183 = io_axi_b_valid ? _GEN_2055 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2184 = io_axi_b_valid ? _GEN_2056 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2185 = io_axi_b_valid ? _GEN_2057 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2186 = io_axi_b_valid ? _GEN_2058 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2187 = io_axi_b_valid ? _GEN_2059 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2188 = io_axi_b_valid ? _GEN_2060 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2189 = io_axi_b_valid ? _GEN_2061 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2190 = io_axi_b_valid ? _GEN_2062 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2191 = io_axi_b_valid ? _GEN_2063 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2192 = io_axi_b_valid ? _GEN_2064 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2193 = io_axi_b_valid ? _GEN_2065 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2194 = io_axi_b_valid ? _GEN_2066 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2195 = io_axi_b_valid ? _GEN_2067 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2196 = io_axi_b_valid ? _GEN_2068 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2197 = io_axi_b_valid ? _GEN_2069 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2198 = io_axi_b_valid ? _GEN_2070 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2199 = io_axi_b_valid ? _GEN_2071 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2200 = io_axi_b_valid ? _GEN_2072 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2201 = io_axi_b_valid ? _GEN_2073 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2202 = io_axi_b_valid ? _GEN_2074 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2203 = io_axi_b_valid ? _GEN_2075 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2204 = io_axi_b_valid ? _GEN_2076 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2205 = io_axi_b_valid ? _GEN_2077 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2206 = io_axi_b_valid ? _GEN_2078 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2207 = io_axi_b_valid ? _GEN_2079 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2208 = io_axi_b_valid ? _GEN_2080 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2209 = io_axi_b_valid ? _GEN_2081 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2210 = io_axi_b_valid ? _GEN_2082 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 406:30]
  wire  _GEN_2211 = io_axi_b_valid ? 1'h0 : fence; // @[playground/src/cache/DCache.scala 145:22 406:30 410:41]
  wire [19:0] _aw_addr_T_1 = _GEN_6610 ? tagRam_0_io_rdata : tagRam_1_io_rdata; // @[playground/src/cache/DCache.scala 418:16]
  wire [31:0] _aw_addr_T_2 = {_aw_addr_T_1,dirty_index,6'h0}; // @[playground/src/cache/DCache.scala 417:25]
  wire [63:0] _GEN_2213 = _GEN_1929 ? data_0_1 : data_0_0; // @[playground/src/cache/DCache.scala 425:{24,24}]
  wire  _GEN_2214 = readsram ? 1'h0 : 1'h1; // @[playground/src/cache/DCache.scala 413:18 414:24 416:20]
  wire [63:0] _GEN_2215 = readsram ? {{32'd0}, _aw_addr_T_2} : _GEN_295; // @[playground/src/cache/DCache.scala 414:24 417:19]
  wire [7:0] _GEN_2216 = readsram ? 8'h7 : _GEN_299; // @[playground/src/cache/DCache.scala 414:24 422:24]
  wire [2:0] _GEN_2217 = readsram ? 3'h3 : _GEN_296; // @[playground/src/cache/DCache.scala 414:24 423:24]
  wire  _GEN_2218 = readsram | _GEN_290; // @[playground/src/cache/DCache.scala 414:24 424:24]
  wire [63:0] _GEN_2219 = readsram ? _GEN_2213 : _GEN_297; // @[playground/src/cache/DCache.scala 414:24 425:24]
  wire [7:0] _GEN_2220 = readsram ? 8'hff : _GEN_298; // @[playground/src/cache/DCache.scala 414:24 426:24]
  wire  _GEN_2221 = readsram ? 1'h0 : _GEN_292; // @[playground/src/cache/DCache.scala 414:24 427:24]
  wire  _GEN_2222 = readsram | _GEN_291; // @[playground/src/cache/DCache.scala 414:24 428:24]
  wire [2:0] _GEN_2223 = readsram ? 3'h0 : bank_wbindex; // @[playground/src/cache/DCache.scala 414:24 429:24 165:29]
  wire  _GEN_2224 = readsram | fence; // @[playground/src/cache/DCache.scala 145:22 414:24 430:24]
  wire  _GEN_2225 = _T_14 ? _GEN_2214 : readsram; // @[playground/src/cache/DCache.scala 148:25 412:36]
  wire [63:0] _GEN_2226 = _T_14 ? _GEN_2215 : _GEN_295; // @[playground/src/cache/DCache.scala 412:36]
  wire [7:0] _GEN_2227 = _T_14 ? _GEN_2216 : _GEN_299; // @[playground/src/cache/DCache.scala 412:36]
  wire [2:0] _GEN_2228 = _T_14 ? _GEN_2217 : _GEN_296; // @[playground/src/cache/DCache.scala 412:36]
  wire  _GEN_2229 = _T_14 ? _GEN_2218 : _GEN_290; // @[playground/src/cache/DCache.scala 412:36]
  wire [63:0] _GEN_2230 = _T_14 ? _GEN_2219 : _GEN_297; // @[playground/src/cache/DCache.scala 412:36]
  wire [7:0] _GEN_2231 = _T_14 ? _GEN_2220 : _GEN_298; // @[playground/src/cache/DCache.scala 412:36]
  wire  _GEN_2232 = _T_14 ? _GEN_2221 : _GEN_292; // @[playground/src/cache/DCache.scala 412:36]
  wire  _GEN_2233 = _T_14 ? _GEN_2222 : _GEN_291; // @[playground/src/cache/DCache.scala 412:36]
  wire [2:0] _GEN_2234 = _T_14 ? _GEN_2223 : bank_wbindex; // @[playground/src/cache/DCache.scala 165:29 412:36]
  wire  _GEN_2235 = _T_14 ? _GEN_2224 : fence; // @[playground/src/cache/DCache.scala 145:22 412:36]
  wire [2:0] _GEN_2236 = _T_14 ? state : 3'h4; // @[playground/src/cache/DCache.scala 412:36 433:15 90:94]
  wire  _GEN_2237 = fence ? _GEN_1865 : _GEN_2229; // @[playground/src/cache/DCache.scala 391:19]
  wire  _GEN_2238 = fence ? _GEN_1951 : _GEN_2233; // @[playground/src/cache/DCache.scala 391:19]
  wire [2:0] _GEN_2239 = fence ? _GEN_1952 : _GEN_2234; // @[playground/src/cache/DCache.scala 391:19]
  wire [63:0] _GEN_2240 = fence ? _GEN_1953 : _GEN_2230; // @[playground/src/cache/DCache.scala 391:19]
  wire  _GEN_2241 = fence ? _GEN_1954 : _GEN_2232; // @[playground/src/cache/DCache.scala 391:19]
  wire  _GEN_2242 = fence ? _GEN_2083 : dirty_0_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2243 = fence ? _GEN_2084 : dirty_0_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2244 = fence ? _GEN_2085 : dirty_1_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2245 = fence ? _GEN_2086 : dirty_1_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2246 = fence ? _GEN_2087 : dirty_2_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2247 = fence ? _GEN_2088 : dirty_2_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2248 = fence ? _GEN_2089 : dirty_3_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2249 = fence ? _GEN_2090 : dirty_3_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2250 = fence ? _GEN_2091 : dirty_4_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2251 = fence ? _GEN_2092 : dirty_4_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2252 = fence ? _GEN_2093 : dirty_5_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2253 = fence ? _GEN_2094 : dirty_5_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2254 = fence ? _GEN_2095 : dirty_6_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2255 = fence ? _GEN_2096 : dirty_6_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2256 = fence ? _GEN_2097 : dirty_7_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2257 = fence ? _GEN_2098 : dirty_7_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2258 = fence ? _GEN_2099 : dirty_8_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2259 = fence ? _GEN_2100 : dirty_8_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2260 = fence ? _GEN_2101 : dirty_9_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2261 = fence ? _GEN_2102 : dirty_9_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2262 = fence ? _GEN_2103 : dirty_10_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2263 = fence ? _GEN_2104 : dirty_10_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2264 = fence ? _GEN_2105 : dirty_11_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2265 = fence ? _GEN_2106 : dirty_11_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2266 = fence ? _GEN_2107 : dirty_12_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2267 = fence ? _GEN_2108 : dirty_12_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2268 = fence ? _GEN_2109 : dirty_13_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2269 = fence ? _GEN_2110 : dirty_13_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2270 = fence ? _GEN_2111 : dirty_14_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2271 = fence ? _GEN_2112 : dirty_14_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2272 = fence ? _GEN_2113 : dirty_15_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2273 = fence ? _GEN_2114 : dirty_15_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2274 = fence ? _GEN_2115 : dirty_16_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2275 = fence ? _GEN_2116 : dirty_16_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2276 = fence ? _GEN_2117 : dirty_17_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2277 = fence ? _GEN_2118 : dirty_17_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2278 = fence ? _GEN_2119 : dirty_18_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2279 = fence ? _GEN_2120 : dirty_18_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2280 = fence ? _GEN_2121 : dirty_19_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2281 = fence ? _GEN_2122 : dirty_19_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2282 = fence ? _GEN_2123 : dirty_20_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2283 = fence ? _GEN_2124 : dirty_20_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2284 = fence ? _GEN_2125 : dirty_21_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2285 = fence ? _GEN_2126 : dirty_21_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2286 = fence ? _GEN_2127 : dirty_22_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2287 = fence ? _GEN_2128 : dirty_22_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2288 = fence ? _GEN_2129 : dirty_23_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2289 = fence ? _GEN_2130 : dirty_23_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2290 = fence ? _GEN_2131 : dirty_24_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2291 = fence ? _GEN_2132 : dirty_24_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2292 = fence ? _GEN_2133 : dirty_25_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2293 = fence ? _GEN_2134 : dirty_25_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2294 = fence ? _GEN_2135 : dirty_26_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2295 = fence ? _GEN_2136 : dirty_26_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2296 = fence ? _GEN_2137 : dirty_27_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2297 = fence ? _GEN_2138 : dirty_27_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2298 = fence ? _GEN_2139 : dirty_28_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2299 = fence ? _GEN_2140 : dirty_28_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2300 = fence ? _GEN_2141 : dirty_29_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2301 = fence ? _GEN_2142 : dirty_29_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2302 = fence ? _GEN_2143 : dirty_30_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2303 = fence ? _GEN_2144 : dirty_30_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2304 = fence ? _GEN_2145 : dirty_31_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2305 = fence ? _GEN_2146 : dirty_31_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2306 = fence ? _GEN_2147 : dirty_32_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2307 = fence ? _GEN_2148 : dirty_32_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2308 = fence ? _GEN_2149 : dirty_33_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2309 = fence ? _GEN_2150 : dirty_33_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2310 = fence ? _GEN_2151 : dirty_34_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2311 = fence ? _GEN_2152 : dirty_34_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2312 = fence ? _GEN_2153 : dirty_35_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2313 = fence ? _GEN_2154 : dirty_35_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2314 = fence ? _GEN_2155 : dirty_36_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2315 = fence ? _GEN_2156 : dirty_36_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2316 = fence ? _GEN_2157 : dirty_37_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2317 = fence ? _GEN_2158 : dirty_37_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2318 = fence ? _GEN_2159 : dirty_38_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2319 = fence ? _GEN_2160 : dirty_38_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2320 = fence ? _GEN_2161 : dirty_39_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2321 = fence ? _GEN_2162 : dirty_39_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2322 = fence ? _GEN_2163 : dirty_40_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2323 = fence ? _GEN_2164 : dirty_40_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2324 = fence ? _GEN_2165 : dirty_41_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2325 = fence ? _GEN_2166 : dirty_41_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2326 = fence ? _GEN_2167 : dirty_42_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2327 = fence ? _GEN_2168 : dirty_42_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2328 = fence ? _GEN_2169 : dirty_43_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2329 = fence ? _GEN_2170 : dirty_43_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2330 = fence ? _GEN_2171 : dirty_44_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2331 = fence ? _GEN_2172 : dirty_44_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2332 = fence ? _GEN_2173 : dirty_45_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2333 = fence ? _GEN_2174 : dirty_45_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2334 = fence ? _GEN_2175 : dirty_46_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2335 = fence ? _GEN_2176 : dirty_46_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2336 = fence ? _GEN_2177 : dirty_47_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2337 = fence ? _GEN_2178 : dirty_47_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2338 = fence ? _GEN_2179 : dirty_48_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2339 = fence ? _GEN_2180 : dirty_48_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2340 = fence ? _GEN_2181 : dirty_49_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2341 = fence ? _GEN_2182 : dirty_49_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2342 = fence ? _GEN_2183 : dirty_50_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2343 = fence ? _GEN_2184 : dirty_50_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2344 = fence ? _GEN_2185 : dirty_51_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2345 = fence ? _GEN_2186 : dirty_51_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2346 = fence ? _GEN_2187 : dirty_52_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2347 = fence ? _GEN_2188 : dirty_52_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2348 = fence ? _GEN_2189 : dirty_53_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2349 = fence ? _GEN_2190 : dirty_53_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2350 = fence ? _GEN_2191 : dirty_54_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2351 = fence ? _GEN_2192 : dirty_54_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2352 = fence ? _GEN_2193 : dirty_55_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2353 = fence ? _GEN_2194 : dirty_55_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2354 = fence ? _GEN_2195 : dirty_56_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2355 = fence ? _GEN_2196 : dirty_56_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2356 = fence ? _GEN_2197 : dirty_57_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2357 = fence ? _GEN_2198 : dirty_57_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2358 = fence ? _GEN_2199 : dirty_58_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2359 = fence ? _GEN_2200 : dirty_58_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2360 = fence ? _GEN_2201 : dirty_59_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2361 = fence ? _GEN_2202 : dirty_59_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2362 = fence ? _GEN_2203 : dirty_60_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2363 = fence ? _GEN_2204 : dirty_60_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2364 = fence ? _GEN_2205 : dirty_61_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2365 = fence ? _GEN_2206 : dirty_61_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2366 = fence ? _GEN_2207 : dirty_62_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2367 = fence ? _GEN_2208 : dirty_62_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2368 = fence ? _GEN_2209 : dirty_63_0; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2369 = fence ? _GEN_2210 : dirty_63_1; // @[playground/src/cache/DCache.scala 391:19 135:22]
  wire  _GEN_2370 = fence ? _GEN_2211 : _GEN_2235; // @[playground/src/cache/DCache.scala 391:19]
  wire  _GEN_2371 = fence ? readsram : _GEN_2225; // @[playground/src/cache/DCache.scala 391:19 148:25]
  wire [63:0] _GEN_2372 = fence ? _GEN_295 : _GEN_2226; // @[playground/src/cache/DCache.scala 391:19]
  wire [7:0] _GEN_2373 = fence ? _GEN_299 : _GEN_2227; // @[playground/src/cache/DCache.scala 391:19]
  wire [2:0] _GEN_2374 = fence ? _GEN_296 : _GEN_2228; // @[playground/src/cache/DCache.scala 391:19]
  wire [7:0] _GEN_2375 = fence ? _GEN_298 : _GEN_2231; // @[playground/src/cache/DCache.scala 391:19]
  wire [2:0] _GEN_2376 = fence ? state : _GEN_2236; // @[playground/src/cache/DCache.scala 391:19 90:94]
  wire  _GEN_2378 = 6'h1 == replace_index ? lru_1 : lru_0; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2379 = 6'h2 == replace_index ? lru_2 : _GEN_2378; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2380 = 6'h3 == replace_index ? lru_3 : _GEN_2379; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2381 = 6'h4 == replace_index ? lru_4 : _GEN_2380; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2382 = 6'h5 == replace_index ? lru_5 : _GEN_2381; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2383 = 6'h6 == replace_index ? lru_6 : _GEN_2382; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2384 = 6'h7 == replace_index ? lru_7 : _GEN_2383; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2385 = 6'h8 == replace_index ? lru_8 : _GEN_2384; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2386 = 6'h9 == replace_index ? lru_9 : _GEN_2385; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2387 = 6'ha == replace_index ? lru_10 : _GEN_2386; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2388 = 6'hb == replace_index ? lru_11 : _GEN_2387; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2389 = 6'hc == replace_index ? lru_12 : _GEN_2388; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2390 = 6'hd == replace_index ? lru_13 : _GEN_2389; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2391 = 6'he == replace_index ? lru_14 : _GEN_2390; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2392 = 6'hf == replace_index ? lru_15 : _GEN_2391; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2393 = 6'h10 == replace_index ? lru_16 : _GEN_2392; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2394 = 6'h11 == replace_index ? lru_17 : _GEN_2393; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2395 = 6'h12 == replace_index ? lru_18 : _GEN_2394; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2396 = 6'h13 == replace_index ? lru_19 : _GEN_2395; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2397 = 6'h14 == replace_index ? lru_20 : _GEN_2396; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2398 = 6'h15 == replace_index ? lru_21 : _GEN_2397; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2399 = 6'h16 == replace_index ? lru_22 : _GEN_2398; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2400 = 6'h17 == replace_index ? lru_23 : _GEN_2399; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2401 = 6'h18 == replace_index ? lru_24 : _GEN_2400; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2402 = 6'h19 == replace_index ? lru_25 : _GEN_2401; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2403 = 6'h1a == replace_index ? lru_26 : _GEN_2402; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2404 = 6'h1b == replace_index ? lru_27 : _GEN_2403; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2405 = 6'h1c == replace_index ? lru_28 : _GEN_2404; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2406 = 6'h1d == replace_index ? lru_29 : _GEN_2405; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2407 = 6'h1e == replace_index ? lru_30 : _GEN_2406; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2408 = 6'h1f == replace_index ? lru_31 : _GEN_2407; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2409 = 6'h20 == replace_index ? lru_32 : _GEN_2408; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2410 = 6'h21 == replace_index ? lru_33 : _GEN_2409; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2411 = 6'h22 == replace_index ? lru_34 : _GEN_2410; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2412 = 6'h23 == replace_index ? lru_35 : _GEN_2411; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2413 = 6'h24 == replace_index ? lru_36 : _GEN_2412; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2414 = 6'h25 == replace_index ? lru_37 : _GEN_2413; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2415 = 6'h26 == replace_index ? lru_38 : _GEN_2414; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2416 = 6'h27 == replace_index ? lru_39 : _GEN_2415; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2417 = 6'h28 == replace_index ? lru_40 : _GEN_2416; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2418 = 6'h29 == replace_index ? lru_41 : _GEN_2417; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2419 = 6'h2a == replace_index ? lru_42 : _GEN_2418; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2420 = 6'h2b == replace_index ? lru_43 : _GEN_2419; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2421 = 6'h2c == replace_index ? lru_44 : _GEN_2420; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2422 = 6'h2d == replace_index ? lru_45 : _GEN_2421; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2423 = 6'h2e == replace_index ? lru_46 : _GEN_2422; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2424 = 6'h2f == replace_index ? lru_47 : _GEN_2423; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2425 = 6'h30 == replace_index ? lru_48 : _GEN_2424; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2426 = 6'h31 == replace_index ? lru_49 : _GEN_2425; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2427 = 6'h32 == replace_index ? lru_50 : _GEN_2426; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2428 = 6'h33 == replace_index ? lru_51 : _GEN_2427; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2429 = 6'h34 == replace_index ? lru_52 : _GEN_2428; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2430 = 6'h35 == replace_index ? lru_53 : _GEN_2429; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2431 = 6'h36 == replace_index ? lru_54 : _GEN_2430; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2432 = 6'h37 == replace_index ? lru_55 : _GEN_2431; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2433 = 6'h38 == replace_index ? lru_56 : _GEN_2432; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2434 = 6'h39 == replace_index ? lru_57 : _GEN_2433; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2435 = 6'h3a == replace_index ? lru_58 : _GEN_2434; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2436 = 6'h3b == replace_index ? lru_59 : _GEN_2435; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2437 = 6'h3c == replace_index ? lru_60 : _GEN_2436; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2438 = 6'h3d == replace_index ? lru_61 : _GEN_2437; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2439 = 6'h3e == replace_index ? lru_62 : _GEN_2438; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2440 = 6'h3f == replace_index ? lru_63 : _GEN_2439; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2442 = _GEN_6288 & _GEN_2440 ? dirty_0_1 : dirty_0_0; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_6824 = ~_GEN_2440; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2443 = _GEN_6293 & ~_GEN_2440 ? dirty_1_0 : _GEN_2442; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2444 = _GEN_6293 & _GEN_2440 ? dirty_1_1 : _GEN_2443; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2445 = _GEN_6298 & ~_GEN_2440 ? dirty_2_0 : _GEN_2444; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2446 = _GEN_6298 & _GEN_2440 ? dirty_2_1 : _GEN_2445; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2447 = _GEN_6303 & ~_GEN_2440 ? dirty_3_0 : _GEN_2446; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2448 = _GEN_6303 & _GEN_2440 ? dirty_3_1 : _GEN_2447; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2449 = _GEN_6308 & ~_GEN_2440 ? dirty_4_0 : _GEN_2448; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2450 = _GEN_6308 & _GEN_2440 ? dirty_4_1 : _GEN_2449; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2451 = _GEN_6313 & ~_GEN_2440 ? dirty_5_0 : _GEN_2450; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2452 = _GEN_6313 & _GEN_2440 ? dirty_5_1 : _GEN_2451; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2453 = _GEN_6318 & ~_GEN_2440 ? dirty_6_0 : _GEN_2452; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2454 = _GEN_6318 & _GEN_2440 ? dirty_6_1 : _GEN_2453; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2455 = _GEN_6323 & ~_GEN_2440 ? dirty_7_0 : _GEN_2454; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2456 = _GEN_6323 & _GEN_2440 ? dirty_7_1 : _GEN_2455; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2457 = _GEN_6328 & ~_GEN_2440 ? dirty_8_0 : _GEN_2456; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2458 = _GEN_6328 & _GEN_2440 ? dirty_8_1 : _GEN_2457; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2459 = _GEN_6333 & ~_GEN_2440 ? dirty_9_0 : _GEN_2458; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2460 = _GEN_6333 & _GEN_2440 ? dirty_9_1 : _GEN_2459; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2461 = _GEN_6338 & ~_GEN_2440 ? dirty_10_0 : _GEN_2460; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2462 = _GEN_6338 & _GEN_2440 ? dirty_10_1 : _GEN_2461; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2463 = _GEN_6343 & ~_GEN_2440 ? dirty_11_0 : _GEN_2462; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2464 = _GEN_6343 & _GEN_2440 ? dirty_11_1 : _GEN_2463; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2465 = _GEN_6348 & ~_GEN_2440 ? dirty_12_0 : _GEN_2464; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2466 = _GEN_6348 & _GEN_2440 ? dirty_12_1 : _GEN_2465; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2467 = _GEN_6353 & ~_GEN_2440 ? dirty_13_0 : _GEN_2466; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2468 = _GEN_6353 & _GEN_2440 ? dirty_13_1 : _GEN_2467; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2469 = _GEN_6358 & ~_GEN_2440 ? dirty_14_0 : _GEN_2468; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2470 = _GEN_6358 & _GEN_2440 ? dirty_14_1 : _GEN_2469; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2471 = _GEN_6363 & ~_GEN_2440 ? dirty_15_0 : _GEN_2470; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2472 = _GEN_6363 & _GEN_2440 ? dirty_15_1 : _GEN_2471; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2473 = _GEN_6368 & ~_GEN_2440 ? dirty_16_0 : _GEN_2472; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2474 = _GEN_6368 & _GEN_2440 ? dirty_16_1 : _GEN_2473; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2475 = _GEN_6373 & ~_GEN_2440 ? dirty_17_0 : _GEN_2474; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2476 = _GEN_6373 & _GEN_2440 ? dirty_17_1 : _GEN_2475; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2477 = _GEN_6378 & ~_GEN_2440 ? dirty_18_0 : _GEN_2476; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2478 = _GEN_6378 & _GEN_2440 ? dirty_18_1 : _GEN_2477; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2479 = _GEN_6383 & ~_GEN_2440 ? dirty_19_0 : _GEN_2478; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2480 = _GEN_6383 & _GEN_2440 ? dirty_19_1 : _GEN_2479; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2481 = _GEN_6388 & ~_GEN_2440 ? dirty_20_0 : _GEN_2480; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2482 = _GEN_6388 & _GEN_2440 ? dirty_20_1 : _GEN_2481; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2483 = _GEN_6393 & ~_GEN_2440 ? dirty_21_0 : _GEN_2482; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2484 = _GEN_6393 & _GEN_2440 ? dirty_21_1 : _GEN_2483; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2485 = _GEN_6398 & ~_GEN_2440 ? dirty_22_0 : _GEN_2484; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2486 = _GEN_6398 & _GEN_2440 ? dirty_22_1 : _GEN_2485; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2487 = _GEN_6403 & ~_GEN_2440 ? dirty_23_0 : _GEN_2486; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2488 = _GEN_6403 & _GEN_2440 ? dirty_23_1 : _GEN_2487; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2489 = _GEN_6408 & ~_GEN_2440 ? dirty_24_0 : _GEN_2488; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2490 = _GEN_6408 & _GEN_2440 ? dirty_24_1 : _GEN_2489; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2491 = _GEN_6413 & ~_GEN_2440 ? dirty_25_0 : _GEN_2490; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2492 = _GEN_6413 & _GEN_2440 ? dirty_25_1 : _GEN_2491; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2493 = _GEN_6418 & ~_GEN_2440 ? dirty_26_0 : _GEN_2492; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2494 = _GEN_6418 & _GEN_2440 ? dirty_26_1 : _GEN_2493; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2495 = _GEN_6423 & ~_GEN_2440 ? dirty_27_0 : _GEN_2494; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2496 = _GEN_6423 & _GEN_2440 ? dirty_27_1 : _GEN_2495; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2497 = _GEN_6428 & ~_GEN_2440 ? dirty_28_0 : _GEN_2496; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2498 = _GEN_6428 & _GEN_2440 ? dirty_28_1 : _GEN_2497; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2499 = _GEN_6433 & ~_GEN_2440 ? dirty_29_0 : _GEN_2498; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2500 = _GEN_6433 & _GEN_2440 ? dirty_29_1 : _GEN_2499; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2501 = _GEN_6438 & ~_GEN_2440 ? dirty_30_0 : _GEN_2500; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2502 = _GEN_6438 & _GEN_2440 ? dirty_30_1 : _GEN_2501; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2503 = _GEN_6443 & ~_GEN_2440 ? dirty_31_0 : _GEN_2502; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2504 = _GEN_6443 & _GEN_2440 ? dirty_31_1 : _GEN_2503; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2505 = _GEN_6448 & ~_GEN_2440 ? dirty_32_0 : _GEN_2504; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2506 = _GEN_6448 & _GEN_2440 ? dirty_32_1 : _GEN_2505; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2507 = _GEN_6453 & ~_GEN_2440 ? dirty_33_0 : _GEN_2506; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2508 = _GEN_6453 & _GEN_2440 ? dirty_33_1 : _GEN_2507; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2509 = _GEN_6458 & ~_GEN_2440 ? dirty_34_0 : _GEN_2508; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2510 = _GEN_6458 & _GEN_2440 ? dirty_34_1 : _GEN_2509; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2511 = _GEN_6463 & ~_GEN_2440 ? dirty_35_0 : _GEN_2510; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2512 = _GEN_6463 & _GEN_2440 ? dirty_35_1 : _GEN_2511; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2513 = _GEN_6468 & ~_GEN_2440 ? dirty_36_0 : _GEN_2512; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2514 = _GEN_6468 & _GEN_2440 ? dirty_36_1 : _GEN_2513; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2515 = _GEN_6473 & ~_GEN_2440 ? dirty_37_0 : _GEN_2514; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2516 = _GEN_6473 & _GEN_2440 ? dirty_37_1 : _GEN_2515; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2517 = _GEN_6478 & ~_GEN_2440 ? dirty_38_0 : _GEN_2516; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2518 = _GEN_6478 & _GEN_2440 ? dirty_38_1 : _GEN_2517; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2519 = _GEN_6483 & ~_GEN_2440 ? dirty_39_0 : _GEN_2518; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2520 = _GEN_6483 & _GEN_2440 ? dirty_39_1 : _GEN_2519; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2521 = _GEN_6488 & ~_GEN_2440 ? dirty_40_0 : _GEN_2520; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2522 = _GEN_6488 & _GEN_2440 ? dirty_40_1 : _GEN_2521; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2523 = _GEN_6493 & ~_GEN_2440 ? dirty_41_0 : _GEN_2522; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2524 = _GEN_6493 & _GEN_2440 ? dirty_41_1 : _GEN_2523; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2525 = _GEN_6498 & ~_GEN_2440 ? dirty_42_0 : _GEN_2524; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2526 = _GEN_6498 & _GEN_2440 ? dirty_42_1 : _GEN_2525; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2527 = _GEN_6503 & ~_GEN_2440 ? dirty_43_0 : _GEN_2526; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2528 = _GEN_6503 & _GEN_2440 ? dirty_43_1 : _GEN_2527; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2529 = _GEN_6508 & ~_GEN_2440 ? dirty_44_0 : _GEN_2528; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2530 = _GEN_6508 & _GEN_2440 ? dirty_44_1 : _GEN_2529; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2531 = _GEN_6513 & ~_GEN_2440 ? dirty_45_0 : _GEN_2530; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2532 = _GEN_6513 & _GEN_2440 ? dirty_45_1 : _GEN_2531; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2533 = _GEN_6518 & ~_GEN_2440 ? dirty_46_0 : _GEN_2532; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2534 = _GEN_6518 & _GEN_2440 ? dirty_46_1 : _GEN_2533; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2535 = _GEN_6523 & ~_GEN_2440 ? dirty_47_0 : _GEN_2534; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2536 = _GEN_6523 & _GEN_2440 ? dirty_47_1 : _GEN_2535; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2537 = _GEN_6528 & ~_GEN_2440 ? dirty_48_0 : _GEN_2536; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2538 = _GEN_6528 & _GEN_2440 ? dirty_48_1 : _GEN_2537; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2539 = _GEN_6533 & ~_GEN_2440 ? dirty_49_0 : _GEN_2538; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2540 = _GEN_6533 & _GEN_2440 ? dirty_49_1 : _GEN_2539; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2541 = _GEN_6538 & ~_GEN_2440 ? dirty_50_0 : _GEN_2540; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2542 = _GEN_6538 & _GEN_2440 ? dirty_50_1 : _GEN_2541; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2543 = _GEN_6543 & ~_GEN_2440 ? dirty_51_0 : _GEN_2542; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2544 = _GEN_6543 & _GEN_2440 ? dirty_51_1 : _GEN_2543; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2545 = _GEN_6548 & ~_GEN_2440 ? dirty_52_0 : _GEN_2544; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2546 = _GEN_6548 & _GEN_2440 ? dirty_52_1 : _GEN_2545; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2547 = _GEN_6553 & ~_GEN_2440 ? dirty_53_0 : _GEN_2546; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2548 = _GEN_6553 & _GEN_2440 ? dirty_53_1 : _GEN_2547; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2549 = _GEN_6558 & ~_GEN_2440 ? dirty_54_0 : _GEN_2548; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2550 = _GEN_6558 & _GEN_2440 ? dirty_54_1 : _GEN_2549; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2551 = _GEN_6563 & ~_GEN_2440 ? dirty_55_0 : _GEN_2550; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2552 = _GEN_6563 & _GEN_2440 ? dirty_55_1 : _GEN_2551; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2553 = _GEN_6568 & ~_GEN_2440 ? dirty_56_0 : _GEN_2552; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2554 = _GEN_6568 & _GEN_2440 ? dirty_56_1 : _GEN_2553; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2555 = _GEN_6573 & ~_GEN_2440 ? dirty_57_0 : _GEN_2554; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2556 = _GEN_6573 & _GEN_2440 ? dirty_57_1 : _GEN_2555; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2557 = _GEN_6578 & ~_GEN_2440 ? dirty_58_0 : _GEN_2556; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2558 = _GEN_6578 & _GEN_2440 ? dirty_58_1 : _GEN_2557; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2559 = _GEN_6583 & ~_GEN_2440 ? dirty_59_0 : _GEN_2558; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2560 = _GEN_6583 & _GEN_2440 ? dirty_59_1 : _GEN_2559; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2561 = _GEN_6588 & ~_GEN_2440 ? dirty_60_0 : _GEN_2560; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2562 = _GEN_6588 & _GEN_2440 ? dirty_60_1 : _GEN_2561; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2563 = _GEN_6593 & ~_GEN_2440 ? dirty_61_0 : _GEN_2562; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2564 = _GEN_6593 & _GEN_2440 ? dirty_61_1 : _GEN_2563; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2565 = _GEN_6598 & ~_GEN_2440 ? dirty_62_0 : _GEN_2564; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2566 = _GEN_6598 & _GEN_2440 ? dirty_62_1 : _GEN_2565; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2567 = _GEN_6603 & ~_GEN_2440 ? dirty_63_0 : _GEN_2566; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire  _GEN_2568 = _GEN_6603 & _GEN_2440 ? dirty_63_1 : _GEN_2567; // @[playground/src/cache/DCache.scala 440:{31,31}]
  wire [63:0] _GEN_2571 = 3'h1 == _bank_wbindex_T_1 ? bank_wbdata_1 : bank_wbdata_0; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2572 = 3'h2 == _bank_wbindex_T_1 ? bank_wbdata_2 : _GEN_2571; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2573 = 3'h3 == _bank_wbindex_T_1 ? bank_wbdata_3 : _GEN_2572; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2574 = 3'h4 == _bank_wbindex_T_1 ? bank_wbdata_4 : _GEN_2573; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2575 = 3'h5 == _bank_wbindex_T_1 ? bank_wbdata_5 : _GEN_2574; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2576 = 3'h6 == _bank_wbindex_T_1 ? bank_wbdata_6 : _GEN_2575; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2577 = 3'h7 == _bank_wbindex_T_1 ? bank_wbdata_7 : _GEN_2576; // @[playground/src/cache/DCache.scala 449:{30,30}]
  wire [63:0] _GEN_2580 = w_last ? _GEN_297 : _GEN_2577; // @[playground/src/cache/DCache.scala 445:28 449:30]
  wire [63:0] _GEN_2584 = _T_1 ? _GEN_2580 : _GEN_297; // @[playground/src/cache/DCache.scala 444:33]
  wire  _GEN_2586 = _GEN_6288 & _GEN_6824 ? 1'h0 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2587 = _GEN_6288 & _GEN_2440 ? 1'h0 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2588 = _GEN_6293 & _GEN_6824 ? 1'h0 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2589 = _GEN_6293 & _GEN_2440 ? 1'h0 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2590 = _GEN_6298 & _GEN_6824 ? 1'h0 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2591 = _GEN_6298 & _GEN_2440 ? 1'h0 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2592 = _GEN_6303 & _GEN_6824 ? 1'h0 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2593 = _GEN_6303 & _GEN_2440 ? 1'h0 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2594 = _GEN_6308 & _GEN_6824 ? 1'h0 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2595 = _GEN_6308 & _GEN_2440 ? 1'h0 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2596 = _GEN_6313 & _GEN_6824 ? 1'h0 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2597 = _GEN_6313 & _GEN_2440 ? 1'h0 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2598 = _GEN_6318 & _GEN_6824 ? 1'h0 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2599 = _GEN_6318 & _GEN_2440 ? 1'h0 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2600 = _GEN_6323 & _GEN_6824 ? 1'h0 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2601 = _GEN_6323 & _GEN_2440 ? 1'h0 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2602 = _GEN_6328 & _GEN_6824 ? 1'h0 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2603 = _GEN_6328 & _GEN_2440 ? 1'h0 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2604 = _GEN_6333 & _GEN_6824 ? 1'h0 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2605 = _GEN_6333 & _GEN_2440 ? 1'h0 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2606 = _GEN_6338 & _GEN_6824 ? 1'h0 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2607 = _GEN_6338 & _GEN_2440 ? 1'h0 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2608 = _GEN_6343 & _GEN_6824 ? 1'h0 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2609 = _GEN_6343 & _GEN_2440 ? 1'h0 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2610 = _GEN_6348 & _GEN_6824 ? 1'h0 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2611 = _GEN_6348 & _GEN_2440 ? 1'h0 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2612 = _GEN_6353 & _GEN_6824 ? 1'h0 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2613 = _GEN_6353 & _GEN_2440 ? 1'h0 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2614 = _GEN_6358 & _GEN_6824 ? 1'h0 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2615 = _GEN_6358 & _GEN_2440 ? 1'h0 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2616 = _GEN_6363 & _GEN_6824 ? 1'h0 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2617 = _GEN_6363 & _GEN_2440 ? 1'h0 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2618 = _GEN_6368 & _GEN_6824 ? 1'h0 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2619 = _GEN_6368 & _GEN_2440 ? 1'h0 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2620 = _GEN_6373 & _GEN_6824 ? 1'h0 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2621 = _GEN_6373 & _GEN_2440 ? 1'h0 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2622 = _GEN_6378 & _GEN_6824 ? 1'h0 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2623 = _GEN_6378 & _GEN_2440 ? 1'h0 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2624 = _GEN_6383 & _GEN_6824 ? 1'h0 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2625 = _GEN_6383 & _GEN_2440 ? 1'h0 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2626 = _GEN_6388 & _GEN_6824 ? 1'h0 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2627 = _GEN_6388 & _GEN_2440 ? 1'h0 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2628 = _GEN_6393 & _GEN_6824 ? 1'h0 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2629 = _GEN_6393 & _GEN_2440 ? 1'h0 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2630 = _GEN_6398 & _GEN_6824 ? 1'h0 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2631 = _GEN_6398 & _GEN_2440 ? 1'h0 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2632 = _GEN_6403 & _GEN_6824 ? 1'h0 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2633 = _GEN_6403 & _GEN_2440 ? 1'h0 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2634 = _GEN_6408 & _GEN_6824 ? 1'h0 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2635 = _GEN_6408 & _GEN_2440 ? 1'h0 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2636 = _GEN_6413 & _GEN_6824 ? 1'h0 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2637 = _GEN_6413 & _GEN_2440 ? 1'h0 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2638 = _GEN_6418 & _GEN_6824 ? 1'h0 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2639 = _GEN_6418 & _GEN_2440 ? 1'h0 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2640 = _GEN_6423 & _GEN_6824 ? 1'h0 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2641 = _GEN_6423 & _GEN_2440 ? 1'h0 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2642 = _GEN_6428 & _GEN_6824 ? 1'h0 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2643 = _GEN_6428 & _GEN_2440 ? 1'h0 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2644 = _GEN_6433 & _GEN_6824 ? 1'h0 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2645 = _GEN_6433 & _GEN_2440 ? 1'h0 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2646 = _GEN_6438 & _GEN_6824 ? 1'h0 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2647 = _GEN_6438 & _GEN_2440 ? 1'h0 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2648 = _GEN_6443 & _GEN_6824 ? 1'h0 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2649 = _GEN_6443 & _GEN_2440 ? 1'h0 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2650 = _GEN_6448 & _GEN_6824 ? 1'h0 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2651 = _GEN_6448 & _GEN_2440 ? 1'h0 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2652 = _GEN_6453 & _GEN_6824 ? 1'h0 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2653 = _GEN_6453 & _GEN_2440 ? 1'h0 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2654 = _GEN_6458 & _GEN_6824 ? 1'h0 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2655 = _GEN_6458 & _GEN_2440 ? 1'h0 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2656 = _GEN_6463 & _GEN_6824 ? 1'h0 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2657 = _GEN_6463 & _GEN_2440 ? 1'h0 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2658 = _GEN_6468 & _GEN_6824 ? 1'h0 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2659 = _GEN_6468 & _GEN_2440 ? 1'h0 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2660 = _GEN_6473 & _GEN_6824 ? 1'h0 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2661 = _GEN_6473 & _GEN_2440 ? 1'h0 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2662 = _GEN_6478 & _GEN_6824 ? 1'h0 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2663 = _GEN_6478 & _GEN_2440 ? 1'h0 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2664 = _GEN_6483 & _GEN_6824 ? 1'h0 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2665 = _GEN_6483 & _GEN_2440 ? 1'h0 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2666 = _GEN_6488 & _GEN_6824 ? 1'h0 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2667 = _GEN_6488 & _GEN_2440 ? 1'h0 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2668 = _GEN_6493 & _GEN_6824 ? 1'h0 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2669 = _GEN_6493 & _GEN_2440 ? 1'h0 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2670 = _GEN_6498 & _GEN_6824 ? 1'h0 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2671 = _GEN_6498 & _GEN_2440 ? 1'h0 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2672 = _GEN_6503 & _GEN_6824 ? 1'h0 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2673 = _GEN_6503 & _GEN_2440 ? 1'h0 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2674 = _GEN_6508 & _GEN_6824 ? 1'h0 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2675 = _GEN_6508 & _GEN_2440 ? 1'h0 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2676 = _GEN_6513 & _GEN_6824 ? 1'h0 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2677 = _GEN_6513 & _GEN_2440 ? 1'h0 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2678 = _GEN_6518 & _GEN_6824 ? 1'h0 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2679 = _GEN_6518 & _GEN_2440 ? 1'h0 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2680 = _GEN_6523 & _GEN_6824 ? 1'h0 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2681 = _GEN_6523 & _GEN_2440 ? 1'h0 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2682 = _GEN_6528 & _GEN_6824 ? 1'h0 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2683 = _GEN_6528 & _GEN_2440 ? 1'h0 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2684 = _GEN_6533 & _GEN_6824 ? 1'h0 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2685 = _GEN_6533 & _GEN_2440 ? 1'h0 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2686 = _GEN_6538 & _GEN_6824 ? 1'h0 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2687 = _GEN_6538 & _GEN_2440 ? 1'h0 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2688 = _GEN_6543 & _GEN_6824 ? 1'h0 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2689 = _GEN_6543 & _GEN_2440 ? 1'h0 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2690 = _GEN_6548 & _GEN_6824 ? 1'h0 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2691 = _GEN_6548 & _GEN_2440 ? 1'h0 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2692 = _GEN_6553 & _GEN_6824 ? 1'h0 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2693 = _GEN_6553 & _GEN_2440 ? 1'h0 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2694 = _GEN_6558 & _GEN_6824 ? 1'h0 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2695 = _GEN_6558 & _GEN_2440 ? 1'h0 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2696 = _GEN_6563 & _GEN_6824 ? 1'h0 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2697 = _GEN_6563 & _GEN_2440 ? 1'h0 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2698 = _GEN_6568 & _GEN_6824 ? 1'h0 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2699 = _GEN_6568 & _GEN_2440 ? 1'h0 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2700 = _GEN_6573 & _GEN_6824 ? 1'h0 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2701 = _GEN_6573 & _GEN_2440 ? 1'h0 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2702 = _GEN_6578 & _GEN_6824 ? 1'h0 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2703 = _GEN_6578 & _GEN_2440 ? 1'h0 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2704 = _GEN_6583 & _GEN_6824 ? 1'h0 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2705 = _GEN_6583 & _GEN_2440 ? 1'h0 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2706 = _GEN_6588 & _GEN_6824 ? 1'h0 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2707 = _GEN_6588 & _GEN_2440 ? 1'h0 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2708 = _GEN_6593 & _GEN_6824 ? 1'h0 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2709 = _GEN_6593 & _GEN_2440 ? 1'h0 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2710 = _GEN_6598 & _GEN_6824 ? 1'h0 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2711 = _GEN_6598 & _GEN_2440 ? 1'h0 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2712 = _GEN_6603 & _GEN_6824 ? 1'h0 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2713 = _GEN_6603 & _GEN_2440 ? 1'h0 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 458:{29,29}]
  wire  _GEN_2714 = io_axi_b_valid ? _GEN_2586 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2715 = io_axi_b_valid ? _GEN_2587 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2716 = io_axi_b_valid ? _GEN_2588 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2717 = io_axi_b_valid ? _GEN_2589 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2718 = io_axi_b_valid ? _GEN_2590 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2719 = io_axi_b_valid ? _GEN_2591 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2720 = io_axi_b_valid ? _GEN_2592 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2721 = io_axi_b_valid ? _GEN_2593 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2722 = io_axi_b_valid ? _GEN_2594 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2723 = io_axi_b_valid ? _GEN_2595 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2724 = io_axi_b_valid ? _GEN_2596 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2725 = io_axi_b_valid ? _GEN_2597 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2726 = io_axi_b_valid ? _GEN_2598 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2727 = io_axi_b_valid ? _GEN_2599 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2728 = io_axi_b_valid ? _GEN_2600 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2729 = io_axi_b_valid ? _GEN_2601 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2730 = io_axi_b_valid ? _GEN_2602 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2731 = io_axi_b_valid ? _GEN_2603 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2732 = io_axi_b_valid ? _GEN_2604 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2733 = io_axi_b_valid ? _GEN_2605 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2734 = io_axi_b_valid ? _GEN_2606 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2735 = io_axi_b_valid ? _GEN_2607 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2736 = io_axi_b_valid ? _GEN_2608 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2737 = io_axi_b_valid ? _GEN_2609 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2738 = io_axi_b_valid ? _GEN_2610 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2739 = io_axi_b_valid ? _GEN_2611 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2740 = io_axi_b_valid ? _GEN_2612 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2741 = io_axi_b_valid ? _GEN_2613 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2742 = io_axi_b_valid ? _GEN_2614 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2743 = io_axi_b_valid ? _GEN_2615 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2744 = io_axi_b_valid ? _GEN_2616 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2745 = io_axi_b_valid ? _GEN_2617 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2746 = io_axi_b_valid ? _GEN_2618 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2747 = io_axi_b_valid ? _GEN_2619 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2748 = io_axi_b_valid ? _GEN_2620 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2749 = io_axi_b_valid ? _GEN_2621 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2750 = io_axi_b_valid ? _GEN_2622 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2751 = io_axi_b_valid ? _GEN_2623 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2752 = io_axi_b_valid ? _GEN_2624 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2753 = io_axi_b_valid ? _GEN_2625 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2754 = io_axi_b_valid ? _GEN_2626 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2755 = io_axi_b_valid ? _GEN_2627 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2756 = io_axi_b_valid ? _GEN_2628 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2757 = io_axi_b_valid ? _GEN_2629 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2758 = io_axi_b_valid ? _GEN_2630 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2759 = io_axi_b_valid ? _GEN_2631 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2760 = io_axi_b_valid ? _GEN_2632 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2761 = io_axi_b_valid ? _GEN_2633 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2762 = io_axi_b_valid ? _GEN_2634 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2763 = io_axi_b_valid ? _GEN_2635 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2764 = io_axi_b_valid ? _GEN_2636 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2765 = io_axi_b_valid ? _GEN_2637 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2766 = io_axi_b_valid ? _GEN_2638 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2767 = io_axi_b_valid ? _GEN_2639 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2768 = io_axi_b_valid ? _GEN_2640 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2769 = io_axi_b_valid ? _GEN_2641 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2770 = io_axi_b_valid ? _GEN_2642 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2771 = io_axi_b_valid ? _GEN_2643 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2772 = io_axi_b_valid ? _GEN_2644 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2773 = io_axi_b_valid ? _GEN_2645 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2774 = io_axi_b_valid ? _GEN_2646 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2775 = io_axi_b_valid ? _GEN_2647 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2776 = io_axi_b_valid ? _GEN_2648 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2777 = io_axi_b_valid ? _GEN_2649 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2778 = io_axi_b_valid ? _GEN_2650 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2779 = io_axi_b_valid ? _GEN_2651 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2780 = io_axi_b_valid ? _GEN_2652 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2781 = io_axi_b_valid ? _GEN_2653 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2782 = io_axi_b_valid ? _GEN_2654 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2783 = io_axi_b_valid ? _GEN_2655 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2784 = io_axi_b_valid ? _GEN_2656 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2785 = io_axi_b_valid ? _GEN_2657 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2786 = io_axi_b_valid ? _GEN_2658 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2787 = io_axi_b_valid ? _GEN_2659 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2788 = io_axi_b_valid ? _GEN_2660 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2789 = io_axi_b_valid ? _GEN_2661 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2790 = io_axi_b_valid ? _GEN_2662 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2791 = io_axi_b_valid ? _GEN_2663 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2792 = io_axi_b_valid ? _GEN_2664 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2793 = io_axi_b_valid ? _GEN_2665 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2794 = io_axi_b_valid ? _GEN_2666 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2795 = io_axi_b_valid ? _GEN_2667 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2796 = io_axi_b_valid ? _GEN_2668 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2797 = io_axi_b_valid ? _GEN_2669 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2798 = io_axi_b_valid ? _GEN_2670 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2799 = io_axi_b_valid ? _GEN_2671 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2800 = io_axi_b_valid ? _GEN_2672 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2801 = io_axi_b_valid ? _GEN_2673 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2802 = io_axi_b_valid ? _GEN_2674 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2803 = io_axi_b_valid ? _GEN_2675 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2804 = io_axi_b_valid ? _GEN_2676 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2805 = io_axi_b_valid ? _GEN_2677 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2806 = io_axi_b_valid ? _GEN_2678 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2807 = io_axi_b_valid ? _GEN_2679 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2808 = io_axi_b_valid ? _GEN_2680 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2809 = io_axi_b_valid ? _GEN_2681 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2810 = io_axi_b_valid ? _GEN_2682 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2811 = io_axi_b_valid ? _GEN_2683 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2812 = io_axi_b_valid ? _GEN_2684 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2813 = io_axi_b_valid ? _GEN_2685 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2814 = io_axi_b_valid ? _GEN_2686 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2815 = io_axi_b_valid ? _GEN_2687 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2816 = io_axi_b_valid ? _GEN_2688 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2817 = io_axi_b_valid ? _GEN_2689 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2818 = io_axi_b_valid ? _GEN_2690 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2819 = io_axi_b_valid ? _GEN_2691 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2820 = io_axi_b_valid ? _GEN_2692 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2821 = io_axi_b_valid ? _GEN_2693 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2822 = io_axi_b_valid ? _GEN_2694 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2823 = io_axi_b_valid ? _GEN_2695 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2824 = io_axi_b_valid ? _GEN_2696 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2825 = io_axi_b_valid ? _GEN_2697 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2826 = io_axi_b_valid ? _GEN_2698 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2827 = io_axi_b_valid ? _GEN_2699 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2828 = io_axi_b_valid ? _GEN_2700 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2829 = io_axi_b_valid ? _GEN_2701 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2830 = io_axi_b_valid ? _GEN_2702 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2831 = io_axi_b_valid ? _GEN_2703 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2832 = io_axi_b_valid ? _GEN_2704 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2833 = io_axi_b_valid ? _GEN_2705 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2834 = io_axi_b_valid ? _GEN_2706 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2835 = io_axi_b_valid ? _GEN_2707 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2836 = io_axi_b_valid ? _GEN_2708 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2837 = io_axi_b_valid ? _GEN_2709 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2838 = io_axi_b_valid ? _GEN_2710 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2839 = io_axi_b_valid ? _GEN_2711 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2840 = io_axi_b_valid ? _GEN_2712 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2841 = io_axi_b_valid ? _GEN_2713 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 455:34]
  wire  _GEN_2842 = _GEN_2568 ? _GEN_1865 : _GEN_290; // @[playground/src/cache/DCache.scala 440:31]
  wire  _GEN_2843 = _GEN_2568 ? _GEN_1951 : _GEN_291; // @[playground/src/cache/DCache.scala 440:31]
  wire [2:0] _GEN_2844 = _GEN_2568 ? _GEN_1952 : bank_wbindex; // @[playground/src/cache/DCache.scala 165:29 440:31]
  wire [63:0] _GEN_2845 = _GEN_2568 ? _GEN_2584 : _GEN_297; // @[playground/src/cache/DCache.scala 440:31]
  wire  _GEN_2846 = _GEN_2568 ? _GEN_1954 : _GEN_292; // @[playground/src/cache/DCache.scala 440:31]
  wire  _GEN_2847 = _GEN_2568 ? _GEN_2714 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2848 = _GEN_2568 ? _GEN_2715 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2849 = _GEN_2568 ? _GEN_2716 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2850 = _GEN_2568 ? _GEN_2717 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2851 = _GEN_2568 ? _GEN_2718 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2852 = _GEN_2568 ? _GEN_2719 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2853 = _GEN_2568 ? _GEN_2720 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2854 = _GEN_2568 ? _GEN_2721 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2855 = _GEN_2568 ? _GEN_2722 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2856 = _GEN_2568 ? _GEN_2723 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2857 = _GEN_2568 ? _GEN_2724 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2858 = _GEN_2568 ? _GEN_2725 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2859 = _GEN_2568 ? _GEN_2726 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2860 = _GEN_2568 ? _GEN_2727 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2861 = _GEN_2568 ? _GEN_2728 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2862 = _GEN_2568 ? _GEN_2729 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2863 = _GEN_2568 ? _GEN_2730 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2864 = _GEN_2568 ? _GEN_2731 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2865 = _GEN_2568 ? _GEN_2732 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2866 = _GEN_2568 ? _GEN_2733 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2867 = _GEN_2568 ? _GEN_2734 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2868 = _GEN_2568 ? _GEN_2735 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2869 = _GEN_2568 ? _GEN_2736 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2870 = _GEN_2568 ? _GEN_2737 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2871 = _GEN_2568 ? _GEN_2738 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2872 = _GEN_2568 ? _GEN_2739 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2873 = _GEN_2568 ? _GEN_2740 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2874 = _GEN_2568 ? _GEN_2741 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2875 = _GEN_2568 ? _GEN_2742 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2876 = _GEN_2568 ? _GEN_2743 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2877 = _GEN_2568 ? _GEN_2744 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2878 = _GEN_2568 ? _GEN_2745 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2879 = _GEN_2568 ? _GEN_2746 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2880 = _GEN_2568 ? _GEN_2747 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2881 = _GEN_2568 ? _GEN_2748 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2882 = _GEN_2568 ? _GEN_2749 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2883 = _GEN_2568 ? _GEN_2750 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2884 = _GEN_2568 ? _GEN_2751 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2885 = _GEN_2568 ? _GEN_2752 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2886 = _GEN_2568 ? _GEN_2753 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2887 = _GEN_2568 ? _GEN_2754 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2888 = _GEN_2568 ? _GEN_2755 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2889 = _GEN_2568 ? _GEN_2756 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2890 = _GEN_2568 ? _GEN_2757 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2891 = _GEN_2568 ? _GEN_2758 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2892 = _GEN_2568 ? _GEN_2759 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2893 = _GEN_2568 ? _GEN_2760 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2894 = _GEN_2568 ? _GEN_2761 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2895 = _GEN_2568 ? _GEN_2762 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2896 = _GEN_2568 ? _GEN_2763 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2897 = _GEN_2568 ? _GEN_2764 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2898 = _GEN_2568 ? _GEN_2765 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2899 = _GEN_2568 ? _GEN_2766 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2900 = _GEN_2568 ? _GEN_2767 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2901 = _GEN_2568 ? _GEN_2768 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2902 = _GEN_2568 ? _GEN_2769 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2903 = _GEN_2568 ? _GEN_2770 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2904 = _GEN_2568 ? _GEN_2771 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2905 = _GEN_2568 ? _GEN_2772 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2906 = _GEN_2568 ? _GEN_2773 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2907 = _GEN_2568 ? _GEN_2774 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2908 = _GEN_2568 ? _GEN_2775 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2909 = _GEN_2568 ? _GEN_2776 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2910 = _GEN_2568 ? _GEN_2777 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2911 = _GEN_2568 ? _GEN_2778 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2912 = _GEN_2568 ? _GEN_2779 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2913 = _GEN_2568 ? _GEN_2780 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2914 = _GEN_2568 ? _GEN_2781 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2915 = _GEN_2568 ? _GEN_2782 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2916 = _GEN_2568 ? _GEN_2783 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2917 = _GEN_2568 ? _GEN_2784 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2918 = _GEN_2568 ? _GEN_2785 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2919 = _GEN_2568 ? _GEN_2786 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2920 = _GEN_2568 ? _GEN_2787 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2921 = _GEN_2568 ? _GEN_2788 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2922 = _GEN_2568 ? _GEN_2789 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2923 = _GEN_2568 ? _GEN_2790 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2924 = _GEN_2568 ? _GEN_2791 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2925 = _GEN_2568 ? _GEN_2792 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2926 = _GEN_2568 ? _GEN_2793 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2927 = _GEN_2568 ? _GEN_2794 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2928 = _GEN_2568 ? _GEN_2795 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2929 = _GEN_2568 ? _GEN_2796 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2930 = _GEN_2568 ? _GEN_2797 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2931 = _GEN_2568 ? _GEN_2798 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2932 = _GEN_2568 ? _GEN_2799 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2933 = _GEN_2568 ? _GEN_2800 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2934 = _GEN_2568 ? _GEN_2801 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2935 = _GEN_2568 ? _GEN_2802 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2936 = _GEN_2568 ? _GEN_2803 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2937 = _GEN_2568 ? _GEN_2804 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2938 = _GEN_2568 ? _GEN_2805 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2939 = _GEN_2568 ? _GEN_2806 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2940 = _GEN_2568 ? _GEN_2807 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2941 = _GEN_2568 ? _GEN_2808 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2942 = _GEN_2568 ? _GEN_2809 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2943 = _GEN_2568 ? _GEN_2810 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2944 = _GEN_2568 ? _GEN_2811 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2945 = _GEN_2568 ? _GEN_2812 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2946 = _GEN_2568 ? _GEN_2813 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2947 = _GEN_2568 ? _GEN_2814 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2948 = _GEN_2568 ? _GEN_2815 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2949 = _GEN_2568 ? _GEN_2816 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2950 = _GEN_2568 ? _GEN_2817 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2951 = _GEN_2568 ? _GEN_2818 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2952 = _GEN_2568 ? _GEN_2819 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2953 = _GEN_2568 ? _GEN_2820 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2954 = _GEN_2568 ? _GEN_2821 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2955 = _GEN_2568 ? _GEN_2822 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2956 = _GEN_2568 ? _GEN_2823 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2957 = _GEN_2568 ? _GEN_2824 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2958 = _GEN_2568 ? _GEN_2825 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2959 = _GEN_2568 ? _GEN_2826 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2960 = _GEN_2568 ? _GEN_2827 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2961 = _GEN_2568 ? _GEN_2828 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2962 = _GEN_2568 ? _GEN_2829 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2963 = _GEN_2568 ? _GEN_2830 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2964 = _GEN_2568 ? _GEN_2831 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2965 = _GEN_2568 ? _GEN_2832 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2966 = _GEN_2568 ? _GEN_2833 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2967 = _GEN_2568 ? _GEN_2834 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2968 = _GEN_2568 ? _GEN_2835 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2969 = _GEN_2568 ? _GEN_2836 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2970 = _GEN_2568 ? _GEN_2837 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2971 = _GEN_2568 ? _GEN_2838 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2972 = _GEN_2568 ? _GEN_2839 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2973 = _GEN_2568 ? _GEN_2840 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _GEN_2974 = _GEN_2568 ? _GEN_2841 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 440:31]
  wire  _T_34 = io_axi_ar_ready & io_axi_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _GEN_2975 = ~_GEN_2440 ? 1'h0 : tag_wstrb_0; // @[playground/src/cache/DCache.scala 182:27 462:{36,36}]
  wire  _GEN_2976 = _GEN_2440 ? 1'h0 : tag_wstrb_1; // @[playground/src/cache/DCache.scala 182:27 462:{36,36}]
  wire  _GEN_2977 = _T_34 ? _GEN_2975 : tag_wstrb_0; // @[playground/src/cache/DCache.scala 182:27 461:32]
  wire  _GEN_2978 = _T_34 ? _GEN_2976 : tag_wstrb_1; // @[playground/src/cache/DCache.scala 182:27 461:32]
  wire  _GEN_2979 = _T_34 ? 1'h0 : arvalid; // @[playground/src/cache/DCache.scala 260:24 461:32 463:36]
  wire [7:0] _GEN_2980 = ~_GEN_2440 ? 8'h0 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22 468:{40,40}]
  wire [7:0] _GEN_2981 = _GEN_2440 ? 8'h0 : burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22 468:{40,40}]
  wire [7:0] _GEN_2983 = _GEN_2440 ? burst_wstrb_1 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 470:{68,68}]
  wire [8:0] _burst_wstrb_T = {_GEN_2983, 1'h0}; // @[playground/src/cache/DCache.scala 470:68]
  wire [7:0] _GEN_2984 = ~_GEN_2440 ? _burst_wstrb_T[7:0] : burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22 470:{40,40}]
  wire [7:0] _GEN_2985 = _GEN_2440 ? _burst_wstrb_T[7:0] : burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22 470:{40,40}]
  wire  _GEN_2986 = io_axi_r_bits_last ? 1'h0 : rready; // @[playground/src/cache/DCache.scala 263:23 466:38 467:40]
  wire [7:0] _GEN_2987 = io_axi_r_bits_last ? _GEN_2980 : _GEN_2984; // @[playground/src/cache/DCache.scala 466:38]
  wire [7:0] _GEN_2988 = io_axi_r_bits_last ? _GEN_2981 : _GEN_2985; // @[playground/src/cache/DCache.scala 466:38]
  wire  _GEN_2989 = _T_18 ? _GEN_2986 : rready; // @[playground/src/cache/DCache.scala 263:23 465:31]
  wire [7:0] _GEN_2990 = _T_18 ? _GEN_2987 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22 465:31]
  wire [7:0] _GEN_2991 = _T_18 ? _GEN_2988 : burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22 465:31]
  wire  _T_40 = io_axi_r_valid & io_axi_r_bits_last | ~rready; // @[playground/src/cache/DCache.scala 475:55]
  wire  _T_41 = (~_GEN_2568 | io_axi_b_valid) & _T_40; // @[playground/src/cache/DCache.scala 474:48]
  wire  _GEN_3120 = _GEN_6288 & _GEN_6824 | valid_0_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3121 = _GEN_6288 & _GEN_2440 | valid_0_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3122 = _GEN_6293 & _GEN_6824 | valid_1_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3123 = _GEN_6293 & _GEN_2440 | valid_1_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3124 = _GEN_6298 & _GEN_6824 | valid_2_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3125 = _GEN_6298 & _GEN_2440 | valid_2_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3126 = _GEN_6303 & _GEN_6824 | valid_3_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3127 = _GEN_6303 & _GEN_2440 | valid_3_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3128 = _GEN_6308 & _GEN_6824 | valid_4_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3129 = _GEN_6308 & _GEN_2440 | valid_4_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3130 = _GEN_6313 & _GEN_6824 | valid_5_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3131 = _GEN_6313 & _GEN_2440 | valid_5_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3132 = _GEN_6318 & _GEN_6824 | valid_6_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3133 = _GEN_6318 & _GEN_2440 | valid_6_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3134 = _GEN_6323 & _GEN_6824 | valid_7_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3135 = _GEN_6323 & _GEN_2440 | valid_7_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3136 = _GEN_6328 & _GEN_6824 | valid_8_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3137 = _GEN_6328 & _GEN_2440 | valid_8_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3138 = _GEN_6333 & _GEN_6824 | valid_9_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3139 = _GEN_6333 & _GEN_2440 | valid_9_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3140 = _GEN_6338 & _GEN_6824 | valid_10_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3141 = _GEN_6338 & _GEN_2440 | valid_10_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3142 = _GEN_6343 & _GEN_6824 | valid_11_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3143 = _GEN_6343 & _GEN_2440 | valid_11_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3144 = _GEN_6348 & _GEN_6824 | valid_12_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3145 = _GEN_6348 & _GEN_2440 | valid_12_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3146 = _GEN_6353 & _GEN_6824 | valid_13_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3147 = _GEN_6353 & _GEN_2440 | valid_13_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3148 = _GEN_6358 & _GEN_6824 | valid_14_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3149 = _GEN_6358 & _GEN_2440 | valid_14_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3150 = _GEN_6363 & _GEN_6824 | valid_15_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3151 = _GEN_6363 & _GEN_2440 | valid_15_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3152 = _GEN_6368 & _GEN_6824 | valid_16_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3153 = _GEN_6368 & _GEN_2440 | valid_16_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3154 = _GEN_6373 & _GEN_6824 | valid_17_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3155 = _GEN_6373 & _GEN_2440 | valid_17_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3156 = _GEN_6378 & _GEN_6824 | valid_18_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3157 = _GEN_6378 & _GEN_2440 | valid_18_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3158 = _GEN_6383 & _GEN_6824 | valid_19_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3159 = _GEN_6383 & _GEN_2440 | valid_19_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3160 = _GEN_6388 & _GEN_6824 | valid_20_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3161 = _GEN_6388 & _GEN_2440 | valid_20_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3162 = _GEN_6393 & _GEN_6824 | valid_21_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3163 = _GEN_6393 & _GEN_2440 | valid_21_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3164 = _GEN_6398 & _GEN_6824 | valid_22_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3165 = _GEN_6398 & _GEN_2440 | valid_22_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3166 = _GEN_6403 & _GEN_6824 | valid_23_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3167 = _GEN_6403 & _GEN_2440 | valid_23_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3168 = _GEN_6408 & _GEN_6824 | valid_24_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3169 = _GEN_6408 & _GEN_2440 | valid_24_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3170 = _GEN_6413 & _GEN_6824 | valid_25_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3171 = _GEN_6413 & _GEN_2440 | valid_25_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3172 = _GEN_6418 & _GEN_6824 | valid_26_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3173 = _GEN_6418 & _GEN_2440 | valid_26_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3174 = _GEN_6423 & _GEN_6824 | valid_27_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3175 = _GEN_6423 & _GEN_2440 | valid_27_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3176 = _GEN_6428 & _GEN_6824 | valid_28_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3177 = _GEN_6428 & _GEN_2440 | valid_28_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3178 = _GEN_6433 & _GEN_6824 | valid_29_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3179 = _GEN_6433 & _GEN_2440 | valid_29_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3180 = _GEN_6438 & _GEN_6824 | valid_30_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3181 = _GEN_6438 & _GEN_2440 | valid_30_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3182 = _GEN_6443 & _GEN_6824 | valid_31_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3183 = _GEN_6443 & _GEN_2440 | valid_31_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3184 = _GEN_6448 & _GEN_6824 | valid_32_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3185 = _GEN_6448 & _GEN_2440 | valid_32_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3186 = _GEN_6453 & _GEN_6824 | valid_33_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3187 = _GEN_6453 & _GEN_2440 | valid_33_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3188 = _GEN_6458 & _GEN_6824 | valid_34_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3189 = _GEN_6458 & _GEN_2440 | valid_34_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3190 = _GEN_6463 & _GEN_6824 | valid_35_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3191 = _GEN_6463 & _GEN_2440 | valid_35_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3192 = _GEN_6468 & _GEN_6824 | valid_36_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3193 = _GEN_6468 & _GEN_2440 | valid_36_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3194 = _GEN_6473 & _GEN_6824 | valid_37_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3195 = _GEN_6473 & _GEN_2440 | valid_37_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3196 = _GEN_6478 & _GEN_6824 | valid_38_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3197 = _GEN_6478 & _GEN_2440 | valid_38_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3198 = _GEN_6483 & _GEN_6824 | valid_39_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3199 = _GEN_6483 & _GEN_2440 | valid_39_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3200 = _GEN_6488 & _GEN_6824 | valid_40_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3201 = _GEN_6488 & _GEN_2440 | valid_40_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3202 = _GEN_6493 & _GEN_6824 | valid_41_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3203 = _GEN_6493 & _GEN_2440 | valid_41_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3204 = _GEN_6498 & _GEN_6824 | valid_42_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3205 = _GEN_6498 & _GEN_2440 | valid_42_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3206 = _GEN_6503 & _GEN_6824 | valid_43_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3207 = _GEN_6503 & _GEN_2440 | valid_43_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3208 = _GEN_6508 & _GEN_6824 | valid_44_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3209 = _GEN_6508 & _GEN_2440 | valid_44_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3210 = _GEN_6513 & _GEN_6824 | valid_45_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3211 = _GEN_6513 & _GEN_2440 | valid_45_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3212 = _GEN_6518 & _GEN_6824 | valid_46_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3213 = _GEN_6518 & _GEN_2440 | valid_46_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3214 = _GEN_6523 & _GEN_6824 | valid_47_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3215 = _GEN_6523 & _GEN_2440 | valid_47_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3216 = _GEN_6528 & _GEN_6824 | valid_48_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3217 = _GEN_6528 & _GEN_2440 | valid_48_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3218 = _GEN_6533 & _GEN_6824 | valid_49_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3219 = _GEN_6533 & _GEN_2440 | valid_49_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3220 = _GEN_6538 & _GEN_6824 | valid_50_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3221 = _GEN_6538 & _GEN_2440 | valid_50_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3222 = _GEN_6543 & _GEN_6824 | valid_51_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3223 = _GEN_6543 & _GEN_2440 | valid_51_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3224 = _GEN_6548 & _GEN_6824 | valid_52_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3225 = _GEN_6548 & _GEN_2440 | valid_52_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3226 = _GEN_6553 & _GEN_6824 | valid_53_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3227 = _GEN_6553 & _GEN_2440 | valid_53_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3228 = _GEN_6558 & _GEN_6824 | valid_54_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3229 = _GEN_6558 & _GEN_2440 | valid_54_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3230 = _GEN_6563 & _GEN_6824 | valid_55_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3231 = _GEN_6563 & _GEN_2440 | valid_55_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3232 = _GEN_6568 & _GEN_6824 | valid_56_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3233 = _GEN_6568 & _GEN_2440 | valid_56_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3234 = _GEN_6573 & _GEN_6824 | valid_57_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3235 = _GEN_6573 & _GEN_2440 | valid_57_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3236 = _GEN_6578 & _GEN_6824 | valid_58_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3237 = _GEN_6578 & _GEN_2440 | valid_58_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3238 = _GEN_6583 & _GEN_6824 | valid_59_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3239 = _GEN_6583 & _GEN_2440 | valid_59_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3240 = _GEN_6588 & _GEN_6824 | valid_60_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3241 = _GEN_6588 & _GEN_2440 | valid_60_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3242 = _GEN_6593 & _GEN_6824 | valid_61_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3243 = _GEN_6593 & _GEN_2440 | valid_61_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3244 = _GEN_6598 & _GEN_6824 | valid_62_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3245 = _GEN_6598 & _GEN_2440 | valid_62_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3246 = _GEN_6603 & _GEN_6824 | valid_63_0; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire  _GEN_3247 = _GEN_6603 & _GEN_2440 | valid_63_1; // @[playground/src/cache/DCache.scala 134:22 477:{47,47}]
  wire [2:0] _GEN_3248 = ptw_scratch_dcache_wait & _T_7 ? 3'h4 : 3'h0; // @[playground/src/cache/DCache.scala 484:80 485:23 488:41]
  wire  _GEN_3249 = ptw_scratch_dcache_wait & _T_7 & ptw_scratch_dcache_wait; // @[playground/src/cache/DCache.scala 101:28 484:80 487:41]
  wire [2:0] _GEN_3250 = ptw_working & io_cpu_tlb_ptw_access_type != 2'h0 ? 3'h5 : _GEN_3248; // @[playground/src/cache/DCache.scala 480:82 482:21]
  wire  _GEN_3251 = ptw_working & io_cpu_tlb_ptw_access_type != 2'h0 ? ptw_scratch_dcache_wait : _GEN_3249; // @[playground/src/cache/DCache.scala 101:28 480:82]
  wire  _GEN_3252 = _T_41 ? _GEN_3120 : valid_0_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3253 = _T_41 ? _GEN_3121 : valid_0_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3254 = _T_41 ? _GEN_3122 : valid_1_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3255 = _T_41 ? _GEN_3123 : valid_1_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3256 = _T_41 ? _GEN_3124 : valid_2_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3257 = _T_41 ? _GEN_3125 : valid_2_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3258 = _T_41 ? _GEN_3126 : valid_3_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3259 = _T_41 ? _GEN_3127 : valid_3_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3260 = _T_41 ? _GEN_3128 : valid_4_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3261 = _T_41 ? _GEN_3129 : valid_4_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3262 = _T_41 ? _GEN_3130 : valid_5_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3263 = _T_41 ? _GEN_3131 : valid_5_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3264 = _T_41 ? _GEN_3132 : valid_6_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3265 = _T_41 ? _GEN_3133 : valid_6_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3266 = _T_41 ? _GEN_3134 : valid_7_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3267 = _T_41 ? _GEN_3135 : valid_7_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3268 = _T_41 ? _GEN_3136 : valid_8_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3269 = _T_41 ? _GEN_3137 : valid_8_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3270 = _T_41 ? _GEN_3138 : valid_9_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3271 = _T_41 ? _GEN_3139 : valid_9_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3272 = _T_41 ? _GEN_3140 : valid_10_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3273 = _T_41 ? _GEN_3141 : valid_10_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3274 = _T_41 ? _GEN_3142 : valid_11_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3275 = _T_41 ? _GEN_3143 : valid_11_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3276 = _T_41 ? _GEN_3144 : valid_12_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3277 = _T_41 ? _GEN_3145 : valid_12_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3278 = _T_41 ? _GEN_3146 : valid_13_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3279 = _T_41 ? _GEN_3147 : valid_13_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3280 = _T_41 ? _GEN_3148 : valid_14_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3281 = _T_41 ? _GEN_3149 : valid_14_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3282 = _T_41 ? _GEN_3150 : valid_15_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3283 = _T_41 ? _GEN_3151 : valid_15_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3284 = _T_41 ? _GEN_3152 : valid_16_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3285 = _T_41 ? _GEN_3153 : valid_16_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3286 = _T_41 ? _GEN_3154 : valid_17_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3287 = _T_41 ? _GEN_3155 : valid_17_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3288 = _T_41 ? _GEN_3156 : valid_18_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3289 = _T_41 ? _GEN_3157 : valid_18_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3290 = _T_41 ? _GEN_3158 : valid_19_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3291 = _T_41 ? _GEN_3159 : valid_19_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3292 = _T_41 ? _GEN_3160 : valid_20_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3293 = _T_41 ? _GEN_3161 : valid_20_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3294 = _T_41 ? _GEN_3162 : valid_21_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3295 = _T_41 ? _GEN_3163 : valid_21_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3296 = _T_41 ? _GEN_3164 : valid_22_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3297 = _T_41 ? _GEN_3165 : valid_22_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3298 = _T_41 ? _GEN_3166 : valid_23_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3299 = _T_41 ? _GEN_3167 : valid_23_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3300 = _T_41 ? _GEN_3168 : valid_24_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3301 = _T_41 ? _GEN_3169 : valid_24_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3302 = _T_41 ? _GEN_3170 : valid_25_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3303 = _T_41 ? _GEN_3171 : valid_25_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3304 = _T_41 ? _GEN_3172 : valid_26_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3305 = _T_41 ? _GEN_3173 : valid_26_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3306 = _T_41 ? _GEN_3174 : valid_27_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3307 = _T_41 ? _GEN_3175 : valid_27_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3308 = _T_41 ? _GEN_3176 : valid_28_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3309 = _T_41 ? _GEN_3177 : valid_28_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3310 = _T_41 ? _GEN_3178 : valid_29_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3311 = _T_41 ? _GEN_3179 : valid_29_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3312 = _T_41 ? _GEN_3180 : valid_30_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3313 = _T_41 ? _GEN_3181 : valid_30_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3314 = _T_41 ? _GEN_3182 : valid_31_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3315 = _T_41 ? _GEN_3183 : valid_31_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3316 = _T_41 ? _GEN_3184 : valid_32_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3317 = _T_41 ? _GEN_3185 : valid_32_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3318 = _T_41 ? _GEN_3186 : valid_33_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3319 = _T_41 ? _GEN_3187 : valid_33_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3320 = _T_41 ? _GEN_3188 : valid_34_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3321 = _T_41 ? _GEN_3189 : valid_34_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3322 = _T_41 ? _GEN_3190 : valid_35_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3323 = _T_41 ? _GEN_3191 : valid_35_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3324 = _T_41 ? _GEN_3192 : valid_36_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3325 = _T_41 ? _GEN_3193 : valid_36_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3326 = _T_41 ? _GEN_3194 : valid_37_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3327 = _T_41 ? _GEN_3195 : valid_37_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3328 = _T_41 ? _GEN_3196 : valid_38_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3329 = _T_41 ? _GEN_3197 : valid_38_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3330 = _T_41 ? _GEN_3198 : valid_39_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3331 = _T_41 ? _GEN_3199 : valid_39_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3332 = _T_41 ? _GEN_3200 : valid_40_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3333 = _T_41 ? _GEN_3201 : valid_40_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3334 = _T_41 ? _GEN_3202 : valid_41_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3335 = _T_41 ? _GEN_3203 : valid_41_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3336 = _T_41 ? _GEN_3204 : valid_42_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3337 = _T_41 ? _GEN_3205 : valid_42_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3338 = _T_41 ? _GEN_3206 : valid_43_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3339 = _T_41 ? _GEN_3207 : valid_43_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3340 = _T_41 ? _GEN_3208 : valid_44_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3341 = _T_41 ? _GEN_3209 : valid_44_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3342 = _T_41 ? _GEN_3210 : valid_45_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3343 = _T_41 ? _GEN_3211 : valid_45_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3344 = _T_41 ? _GEN_3212 : valid_46_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3345 = _T_41 ? _GEN_3213 : valid_46_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3346 = _T_41 ? _GEN_3214 : valid_47_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3347 = _T_41 ? _GEN_3215 : valid_47_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3348 = _T_41 ? _GEN_3216 : valid_48_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3349 = _T_41 ? _GEN_3217 : valid_48_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3350 = _T_41 ? _GEN_3218 : valid_49_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3351 = _T_41 ? _GEN_3219 : valid_49_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3352 = _T_41 ? _GEN_3220 : valid_50_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3353 = _T_41 ? _GEN_3221 : valid_50_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3354 = _T_41 ? _GEN_3222 : valid_51_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3355 = _T_41 ? _GEN_3223 : valid_51_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3356 = _T_41 ? _GEN_3224 : valid_52_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3357 = _T_41 ? _GEN_3225 : valid_52_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3358 = _T_41 ? _GEN_3226 : valid_53_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3359 = _T_41 ? _GEN_3227 : valid_53_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3360 = _T_41 ? _GEN_3228 : valid_54_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3361 = _T_41 ? _GEN_3229 : valid_54_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3362 = _T_41 ? _GEN_3230 : valid_55_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3363 = _T_41 ? _GEN_3231 : valid_55_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3364 = _T_41 ? _GEN_3232 : valid_56_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3365 = _T_41 ? _GEN_3233 : valid_56_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3366 = _T_41 ? _GEN_3234 : valid_57_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3367 = _T_41 ? _GEN_3235 : valid_57_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3368 = _T_41 ? _GEN_3236 : valid_58_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3369 = _T_41 ? _GEN_3237 : valid_58_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3370 = _T_41 ? _GEN_3238 : valid_59_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3371 = _T_41 ? _GEN_3239 : valid_59_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3372 = _T_41 ? _GEN_3240 : valid_60_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3373 = _T_41 ? _GEN_3241 : valid_60_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3374 = _T_41 ? _GEN_3242 : valid_61_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3375 = _T_41 ? _GEN_3243 : valid_61_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3376 = _T_41 ? _GEN_3244 : valid_62_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3377 = _T_41 ? _GEN_3245 : valid_62_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3378 = _T_41 ? _GEN_3246 : valid_63_0; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3379 = _T_41 ? _GEN_3247 : valid_63_1; // @[playground/src/cache/DCache.scala 476:13 134:22]
  wire  _GEN_3380 = _T_41 ? 1'h0 : do_replace; // @[playground/src/cache/DCache.scala 476:13 170:30 478:47]
  wire  _GEN_3381 = _T_41 ? 1'h0 : ptw_scratch_replace; // @[playground/src/cache/DCache.scala 476:13 101:28 479:47]
  wire [2:0] _GEN_3382 = _T_41 ? _GEN_3250 : state; // @[playground/src/cache/DCache.scala 476:13 90:94]
  wire  _GEN_3383 = _T_41 ? _GEN_3251 : ptw_scratch_dcache_wait; // @[playground/src/cache/DCache.scala 476:13 101:28]
  wire [7:0] _GEN_3384 = ~_GEN_2440 ? 8'h1 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22 502:{38,38}]
  wire [7:0] _GEN_3385 = _GEN_2440 ? 8'h1 : burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22 502:{38,38}]
  wire  _GEN_3386 = _GEN_6824 | tag_wstrb_0; // @[playground/src/cache/DCache.scala 182:27 503:{38,38}]
  wire  _GEN_3387 = _GEN_2440 | tag_wstrb_1; // @[playground/src/cache/DCache.scala 182:27 503:{38,38}]
  wire [31:0] _ar_addr_T_1 = {io_cpu_tlb_paddr[31:6],6'h0}; // @[playground/src/cache/DCache.scala 507:31]
  wire [31:0] _ar_addr_T_2 = {ptw_scratch_paddr_tag,ptw_scratch_paddr_index,6'h0}; // @[playground/src/cache/DCache.scala 511:31]
  wire [31:0] _GEN_3388 = _io_cpu_tlb_ptw_vpn_ready_T ? _ar_addr_T_1 : _ar_addr_T_2; // @[playground/src/cache/DCache.scala 504:32 507:25 511:25]
  wire [19:0] _GEN_3389 = _io_cpu_tlb_ptw_vpn_ready_T ? io_cpu_tlb_ptag : ptw_scratch_paddr_tag; // @[playground/src/cache/DCache.scala 504:32 508:25 512:25]
  wire [63:0] _GEN_3519 = _GEN_2440 ? data_0_1 : data_0_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3521 = _GEN_2440 ? data_1_1 : data_1_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3523 = _GEN_2440 ? data_2_1 : data_2_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3525 = _GEN_2440 ? data_3_1 : data_3_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3527 = _GEN_2440 ? data_4_1 : data_4_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3529 = _GEN_2440 ? data_5_1 : data_5_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3531 = _GEN_2440 ? data_6_1 : data_6_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [63:0] _GEN_3533 = _GEN_2440 ? data_7_1 : data_7_0; // @[playground/src/cache/DCache.scala 516:{55,55}]
  wire [19:0] _GEN_3535 = _GEN_2440 ? tag_1 : tag_0; // @[playground/src/cache/DCache.scala 517:{34,34}]
  wire [31:0] _aw_addr_T_3 = {_GEN_3535,replace_index,6'h0}; // @[playground/src/cache/DCache.scala 517:34]
  wire [63:0] _GEN_3538 = _GEN_2568 ? _GEN_3519 : bank_wbdata_0; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3539 = _GEN_2568 ? _GEN_3521 : bank_wbdata_1; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3540 = _GEN_2568 ? _GEN_3523 : bank_wbdata_2; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3541 = _GEN_2568 ? _GEN_3525 : bank_wbdata_3; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3542 = _GEN_2568 ? _GEN_3527 : bank_wbdata_4; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3543 = _GEN_2568 ? _GEN_3529 : bank_wbdata_5; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3544 = _GEN_2568 ? _GEN_3531 : bank_wbdata_6; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3545 = _GEN_2568 ? _GEN_3533 : bank_wbdata_7; // @[playground/src/cache/DCache.scala 166:29 514:33 516:55]
  wire [63:0] _GEN_3546 = _GEN_2568 ? {{32'd0}, _aw_addr_T_3} : _GEN_295; // @[playground/src/cache/DCache.scala 514:33 517:28]
  wire [7:0] _GEN_3547 = _GEN_2568 ? 8'h7 : _GEN_299; // @[playground/src/cache/DCache.scala 514:33 518:28]
  wire [2:0] _GEN_3548 = _GEN_2568 ? 3'h3 : _GEN_296; // @[playground/src/cache/DCache.scala 514:33 519:28]
  wire  _GEN_3549 = _GEN_2568 | _GEN_290; // @[playground/src/cache/DCache.scala 514:33 520:28]
  wire [63:0] _GEN_3550 = _GEN_2568 ? _GEN_3519 : _GEN_297; // @[playground/src/cache/DCache.scala 514:33 521:28]
  wire [7:0] _GEN_3551 = _GEN_2568 ? 8'hff : _GEN_298; // @[playground/src/cache/DCache.scala 514:33 522:28]
  wire  _GEN_3552 = _GEN_2568 ? 1'h0 : _GEN_292; // @[playground/src/cache/DCache.scala 514:33 523:28]
  wire  _GEN_3553 = _GEN_2568 | _GEN_291; // @[playground/src/cache/DCache.scala 514:33 524:28]
  wire [2:0] _GEN_3554 = _GEN_2568 ? 3'h0 : bank_wbindex; // @[playground/src/cache/DCache.scala 514:33 525:28 165:29]
  wire  _GEN_3555 = readsram | do_replace; // @[playground/src/cache/DCache.scala 495:26 170:30 497:38]
  wire [7:0] _GEN_3556 = readsram ? 8'h7 : ar_len; // @[playground/src/cache/DCache.scala 259:24 495:26 498:38]
  wire [2:0] _GEN_3557 = readsram ? 3'h3 : ar_size; // @[playground/src/cache/DCache.scala 259:24 495:26 499:38]
  wire  _GEN_3558 = readsram | arvalid; // @[playground/src/cache/DCache.scala 260:24 495:26 500:38]
  wire  _GEN_3559 = readsram | rready; // @[playground/src/cache/DCache.scala 263:23 495:26 501:38]
  wire [7:0] _GEN_3560 = readsram ? _GEN_3384 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22 495:26]
  wire [7:0] _GEN_3561 = readsram ? _GEN_3385 : burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22 495:26]
  wire  _GEN_3562 = readsram ? _GEN_3386 : tag_wstrb_0; // @[playground/src/cache/DCache.scala 495:26 182:27]
  wire  _GEN_3563 = readsram ? _GEN_3387 : tag_wstrb_1; // @[playground/src/cache/DCache.scala 495:26 182:27]
  wire [31:0] _GEN_3564 = readsram ? _GEN_3388 : ar_addr; // @[playground/src/cache/DCache.scala 259:24 495:26]
  wire [19:0] _GEN_3565 = readsram ? _GEN_3389 : tag_wdata; // @[playground/src/cache/DCache.scala 495:26 183:27]
  wire [63:0] _GEN_3566 = readsram ? _GEN_3538 : bank_wbdata_0; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3567 = readsram ? _GEN_3539 : bank_wbdata_1; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3568 = readsram ? _GEN_3540 : bank_wbdata_2; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3569 = readsram ? _GEN_3541 : bank_wbdata_3; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3570 = readsram ? _GEN_3542 : bank_wbdata_4; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3571 = readsram ? _GEN_3543 : bank_wbdata_5; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3572 = readsram ? _GEN_3544 : bank_wbdata_6; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3573 = readsram ? _GEN_3545 : bank_wbdata_7; // @[playground/src/cache/DCache.scala 495:26 166:29]
  wire [63:0] _GEN_3574 = readsram ? _GEN_3546 : _GEN_295; // @[playground/src/cache/DCache.scala 495:26]
  wire [7:0] _GEN_3575 = readsram ? _GEN_3547 : _GEN_299; // @[playground/src/cache/DCache.scala 495:26]
  wire [2:0] _GEN_3576 = readsram ? _GEN_3548 : _GEN_296; // @[playground/src/cache/DCache.scala 495:26]
  wire  _GEN_3577 = readsram ? _GEN_3549 : _GEN_290; // @[playground/src/cache/DCache.scala 495:26]
  wire [63:0] _GEN_3578 = readsram ? _GEN_3550 : _GEN_297; // @[playground/src/cache/DCache.scala 495:26]
  wire [7:0] _GEN_3579 = readsram ? _GEN_3551 : _GEN_298; // @[playground/src/cache/DCache.scala 495:26]
  wire  _GEN_3580 = readsram ? _GEN_3552 : _GEN_292; // @[playground/src/cache/DCache.scala 495:26]
  wire  _GEN_3581 = readsram ? _GEN_3553 : _GEN_291; // @[playground/src/cache/DCache.scala 495:26]
  wire [2:0] _GEN_3582 = readsram ? _GEN_3554 : bank_wbindex; // @[playground/src/cache/DCache.scala 495:26 165:29]
  wire  _GEN_3583 = do_replace ? _GEN_2842 : _GEN_3577; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3584 = do_replace ? _GEN_2843 : _GEN_3581; // @[playground/src/cache/DCache.scala 439:26]
  wire [2:0] _GEN_3585 = do_replace ? _GEN_2844 : _GEN_3582; // @[playground/src/cache/DCache.scala 439:26]
  wire [63:0] _GEN_3586 = do_replace ? _GEN_2845 : _GEN_3578; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3587 = do_replace ? _GEN_2846 : _GEN_3580; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3588 = do_replace ? _GEN_2847 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3589 = do_replace ? _GEN_2848 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3590 = do_replace ? _GEN_2849 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3591 = do_replace ? _GEN_2850 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3592 = do_replace ? _GEN_2851 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3593 = do_replace ? _GEN_2852 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3594 = do_replace ? _GEN_2853 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3595 = do_replace ? _GEN_2854 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3596 = do_replace ? _GEN_2855 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3597 = do_replace ? _GEN_2856 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3598 = do_replace ? _GEN_2857 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3599 = do_replace ? _GEN_2858 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3600 = do_replace ? _GEN_2859 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3601 = do_replace ? _GEN_2860 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3602 = do_replace ? _GEN_2861 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3603 = do_replace ? _GEN_2862 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3604 = do_replace ? _GEN_2863 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3605 = do_replace ? _GEN_2864 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3606 = do_replace ? _GEN_2865 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3607 = do_replace ? _GEN_2866 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3608 = do_replace ? _GEN_2867 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3609 = do_replace ? _GEN_2868 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3610 = do_replace ? _GEN_2869 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3611 = do_replace ? _GEN_2870 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3612 = do_replace ? _GEN_2871 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3613 = do_replace ? _GEN_2872 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3614 = do_replace ? _GEN_2873 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3615 = do_replace ? _GEN_2874 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3616 = do_replace ? _GEN_2875 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3617 = do_replace ? _GEN_2876 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3618 = do_replace ? _GEN_2877 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3619 = do_replace ? _GEN_2878 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3620 = do_replace ? _GEN_2879 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3621 = do_replace ? _GEN_2880 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3622 = do_replace ? _GEN_2881 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3623 = do_replace ? _GEN_2882 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3624 = do_replace ? _GEN_2883 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3625 = do_replace ? _GEN_2884 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3626 = do_replace ? _GEN_2885 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3627 = do_replace ? _GEN_2886 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3628 = do_replace ? _GEN_2887 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3629 = do_replace ? _GEN_2888 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3630 = do_replace ? _GEN_2889 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3631 = do_replace ? _GEN_2890 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3632 = do_replace ? _GEN_2891 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3633 = do_replace ? _GEN_2892 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3634 = do_replace ? _GEN_2893 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3635 = do_replace ? _GEN_2894 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3636 = do_replace ? _GEN_2895 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3637 = do_replace ? _GEN_2896 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3638 = do_replace ? _GEN_2897 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3639 = do_replace ? _GEN_2898 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3640 = do_replace ? _GEN_2899 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3641 = do_replace ? _GEN_2900 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3642 = do_replace ? _GEN_2901 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3643 = do_replace ? _GEN_2902 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3644 = do_replace ? _GEN_2903 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3645 = do_replace ? _GEN_2904 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3646 = do_replace ? _GEN_2905 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3647 = do_replace ? _GEN_2906 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3648 = do_replace ? _GEN_2907 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3649 = do_replace ? _GEN_2908 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3650 = do_replace ? _GEN_2909 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3651 = do_replace ? _GEN_2910 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3652 = do_replace ? _GEN_2911 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3653 = do_replace ? _GEN_2912 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3654 = do_replace ? _GEN_2913 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3655 = do_replace ? _GEN_2914 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3656 = do_replace ? _GEN_2915 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3657 = do_replace ? _GEN_2916 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3658 = do_replace ? _GEN_2917 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3659 = do_replace ? _GEN_2918 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3660 = do_replace ? _GEN_2919 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3661 = do_replace ? _GEN_2920 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3662 = do_replace ? _GEN_2921 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3663 = do_replace ? _GEN_2922 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3664 = do_replace ? _GEN_2923 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3665 = do_replace ? _GEN_2924 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3666 = do_replace ? _GEN_2925 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3667 = do_replace ? _GEN_2926 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3668 = do_replace ? _GEN_2927 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3669 = do_replace ? _GEN_2928 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3670 = do_replace ? _GEN_2929 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3671 = do_replace ? _GEN_2930 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3672 = do_replace ? _GEN_2931 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3673 = do_replace ? _GEN_2932 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3674 = do_replace ? _GEN_2933 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3675 = do_replace ? _GEN_2934 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3676 = do_replace ? _GEN_2935 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3677 = do_replace ? _GEN_2936 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3678 = do_replace ? _GEN_2937 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3679 = do_replace ? _GEN_2938 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3680 = do_replace ? _GEN_2939 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3681 = do_replace ? _GEN_2940 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3682 = do_replace ? _GEN_2941 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3683 = do_replace ? _GEN_2942 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3684 = do_replace ? _GEN_2943 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3685 = do_replace ? _GEN_2944 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3686 = do_replace ? _GEN_2945 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3687 = do_replace ? _GEN_2946 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3688 = do_replace ? _GEN_2947 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3689 = do_replace ? _GEN_2948 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3690 = do_replace ? _GEN_2949 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3691 = do_replace ? _GEN_2950 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3692 = do_replace ? _GEN_2951 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3693 = do_replace ? _GEN_2952 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3694 = do_replace ? _GEN_2953 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3695 = do_replace ? _GEN_2954 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3696 = do_replace ? _GEN_2955 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3697 = do_replace ? _GEN_2956 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3698 = do_replace ? _GEN_2957 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3699 = do_replace ? _GEN_2958 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3700 = do_replace ? _GEN_2959 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3701 = do_replace ? _GEN_2960 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3702 = do_replace ? _GEN_2961 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3703 = do_replace ? _GEN_2962 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3704 = do_replace ? _GEN_2963 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3705 = do_replace ? _GEN_2964 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3706 = do_replace ? _GEN_2965 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3707 = do_replace ? _GEN_2966 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3708 = do_replace ? _GEN_2967 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3709 = do_replace ? _GEN_2968 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3710 = do_replace ? _GEN_2969 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3711 = do_replace ? _GEN_2970 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3712 = do_replace ? _GEN_2971 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3713 = do_replace ? _GEN_2972 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3714 = do_replace ? _GEN_2973 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3715 = do_replace ? _GEN_2974 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 439:26]
  wire  _GEN_3716 = do_replace ? _GEN_2977 : _GEN_3562; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3717 = do_replace ? _GEN_2978 : _GEN_3563; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3718 = do_replace ? _GEN_2979 : _GEN_3558; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3719 = do_replace ? _GEN_2989 : _GEN_3559; // @[playground/src/cache/DCache.scala 439:26]
  wire [7:0] _GEN_3720 = do_replace ? _GEN_2990 : _GEN_3560; // @[playground/src/cache/DCache.scala 439:26]
  wire [7:0] _GEN_3721 = do_replace ? _GEN_2991 : _GEN_3561; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3722 = do_replace ? _GEN_3252 : valid_0_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3723 = do_replace ? _GEN_3253 : valid_0_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3724 = do_replace ? _GEN_3254 : valid_1_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3725 = do_replace ? _GEN_3255 : valid_1_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3726 = do_replace ? _GEN_3256 : valid_2_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3727 = do_replace ? _GEN_3257 : valid_2_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3728 = do_replace ? _GEN_3258 : valid_3_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3729 = do_replace ? _GEN_3259 : valid_3_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3730 = do_replace ? _GEN_3260 : valid_4_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3731 = do_replace ? _GEN_3261 : valid_4_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3732 = do_replace ? _GEN_3262 : valid_5_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3733 = do_replace ? _GEN_3263 : valid_5_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3734 = do_replace ? _GEN_3264 : valid_6_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3735 = do_replace ? _GEN_3265 : valid_6_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3736 = do_replace ? _GEN_3266 : valid_7_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3737 = do_replace ? _GEN_3267 : valid_7_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3738 = do_replace ? _GEN_3268 : valid_8_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3739 = do_replace ? _GEN_3269 : valid_8_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3740 = do_replace ? _GEN_3270 : valid_9_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3741 = do_replace ? _GEN_3271 : valid_9_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3742 = do_replace ? _GEN_3272 : valid_10_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3743 = do_replace ? _GEN_3273 : valid_10_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3744 = do_replace ? _GEN_3274 : valid_11_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3745 = do_replace ? _GEN_3275 : valid_11_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3746 = do_replace ? _GEN_3276 : valid_12_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3747 = do_replace ? _GEN_3277 : valid_12_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3748 = do_replace ? _GEN_3278 : valid_13_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3749 = do_replace ? _GEN_3279 : valid_13_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3750 = do_replace ? _GEN_3280 : valid_14_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3751 = do_replace ? _GEN_3281 : valid_14_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3752 = do_replace ? _GEN_3282 : valid_15_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3753 = do_replace ? _GEN_3283 : valid_15_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3754 = do_replace ? _GEN_3284 : valid_16_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3755 = do_replace ? _GEN_3285 : valid_16_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3756 = do_replace ? _GEN_3286 : valid_17_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3757 = do_replace ? _GEN_3287 : valid_17_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3758 = do_replace ? _GEN_3288 : valid_18_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3759 = do_replace ? _GEN_3289 : valid_18_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3760 = do_replace ? _GEN_3290 : valid_19_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3761 = do_replace ? _GEN_3291 : valid_19_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3762 = do_replace ? _GEN_3292 : valid_20_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3763 = do_replace ? _GEN_3293 : valid_20_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3764 = do_replace ? _GEN_3294 : valid_21_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3765 = do_replace ? _GEN_3295 : valid_21_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3766 = do_replace ? _GEN_3296 : valid_22_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3767 = do_replace ? _GEN_3297 : valid_22_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3768 = do_replace ? _GEN_3298 : valid_23_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3769 = do_replace ? _GEN_3299 : valid_23_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3770 = do_replace ? _GEN_3300 : valid_24_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3771 = do_replace ? _GEN_3301 : valid_24_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3772 = do_replace ? _GEN_3302 : valid_25_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3773 = do_replace ? _GEN_3303 : valid_25_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3774 = do_replace ? _GEN_3304 : valid_26_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3775 = do_replace ? _GEN_3305 : valid_26_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3776 = do_replace ? _GEN_3306 : valid_27_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3777 = do_replace ? _GEN_3307 : valid_27_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3778 = do_replace ? _GEN_3308 : valid_28_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3779 = do_replace ? _GEN_3309 : valid_28_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3780 = do_replace ? _GEN_3310 : valid_29_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3781 = do_replace ? _GEN_3311 : valid_29_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3782 = do_replace ? _GEN_3312 : valid_30_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3783 = do_replace ? _GEN_3313 : valid_30_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3784 = do_replace ? _GEN_3314 : valid_31_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3785 = do_replace ? _GEN_3315 : valid_31_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3786 = do_replace ? _GEN_3316 : valid_32_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3787 = do_replace ? _GEN_3317 : valid_32_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3788 = do_replace ? _GEN_3318 : valid_33_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3789 = do_replace ? _GEN_3319 : valid_33_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3790 = do_replace ? _GEN_3320 : valid_34_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3791 = do_replace ? _GEN_3321 : valid_34_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3792 = do_replace ? _GEN_3322 : valid_35_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3793 = do_replace ? _GEN_3323 : valid_35_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3794 = do_replace ? _GEN_3324 : valid_36_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3795 = do_replace ? _GEN_3325 : valid_36_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3796 = do_replace ? _GEN_3326 : valid_37_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3797 = do_replace ? _GEN_3327 : valid_37_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3798 = do_replace ? _GEN_3328 : valid_38_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3799 = do_replace ? _GEN_3329 : valid_38_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3800 = do_replace ? _GEN_3330 : valid_39_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3801 = do_replace ? _GEN_3331 : valid_39_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3802 = do_replace ? _GEN_3332 : valid_40_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3803 = do_replace ? _GEN_3333 : valid_40_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3804 = do_replace ? _GEN_3334 : valid_41_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3805 = do_replace ? _GEN_3335 : valid_41_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3806 = do_replace ? _GEN_3336 : valid_42_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3807 = do_replace ? _GEN_3337 : valid_42_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3808 = do_replace ? _GEN_3338 : valid_43_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3809 = do_replace ? _GEN_3339 : valid_43_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3810 = do_replace ? _GEN_3340 : valid_44_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3811 = do_replace ? _GEN_3341 : valid_44_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3812 = do_replace ? _GEN_3342 : valid_45_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3813 = do_replace ? _GEN_3343 : valid_45_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3814 = do_replace ? _GEN_3344 : valid_46_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3815 = do_replace ? _GEN_3345 : valid_46_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3816 = do_replace ? _GEN_3346 : valid_47_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3817 = do_replace ? _GEN_3347 : valid_47_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3818 = do_replace ? _GEN_3348 : valid_48_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3819 = do_replace ? _GEN_3349 : valid_48_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3820 = do_replace ? _GEN_3350 : valid_49_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3821 = do_replace ? _GEN_3351 : valid_49_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3822 = do_replace ? _GEN_3352 : valid_50_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3823 = do_replace ? _GEN_3353 : valid_50_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3824 = do_replace ? _GEN_3354 : valid_51_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3825 = do_replace ? _GEN_3355 : valid_51_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3826 = do_replace ? _GEN_3356 : valid_52_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3827 = do_replace ? _GEN_3357 : valid_52_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3828 = do_replace ? _GEN_3358 : valid_53_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3829 = do_replace ? _GEN_3359 : valid_53_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3830 = do_replace ? _GEN_3360 : valid_54_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3831 = do_replace ? _GEN_3361 : valid_54_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3832 = do_replace ? _GEN_3362 : valid_55_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3833 = do_replace ? _GEN_3363 : valid_55_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3834 = do_replace ? _GEN_3364 : valid_56_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3835 = do_replace ? _GEN_3365 : valid_56_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3836 = do_replace ? _GEN_3366 : valid_57_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3837 = do_replace ? _GEN_3367 : valid_57_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3838 = do_replace ? _GEN_3368 : valid_58_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3839 = do_replace ? _GEN_3369 : valid_58_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3840 = do_replace ? _GEN_3370 : valid_59_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3841 = do_replace ? _GEN_3371 : valid_59_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3842 = do_replace ? _GEN_3372 : valid_60_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3843 = do_replace ? _GEN_3373 : valid_60_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3844 = do_replace ? _GEN_3374 : valid_61_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3845 = do_replace ? _GEN_3375 : valid_61_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3846 = do_replace ? _GEN_3376 : valid_62_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3847 = do_replace ? _GEN_3377 : valid_62_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3848 = do_replace ? _GEN_3378 : valid_63_0; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3849 = do_replace ? _GEN_3379 : valid_63_1; // @[playground/src/cache/DCache.scala 134:22 439:26]
  wire  _GEN_3850 = do_replace ? _GEN_3380 : _GEN_3555; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3851 = do_replace ? _GEN_3381 : ptw_scratch_replace; // @[playground/src/cache/DCache.scala 439:26 101:28]
  wire [2:0] _GEN_3852 = do_replace ? _GEN_3382 : state; // @[playground/src/cache/DCache.scala 439:26 90:94]
  wire  _GEN_3853 = do_replace ? _GEN_3383 : ptw_scratch_dcache_wait; // @[playground/src/cache/DCache.scala 439:26 101:28]
  wire  _GEN_3854 = do_replace ? readsram : _GEN_2214; // @[playground/src/cache/DCache.scala 148:25 439:26]
  wire [7:0] _GEN_3855 = do_replace ? ar_len : _GEN_3556; // @[playground/src/cache/DCache.scala 259:24 439:26]
  wire [2:0] _GEN_3856 = do_replace ? ar_size : _GEN_3557; // @[playground/src/cache/DCache.scala 259:24 439:26]
  wire [31:0] _GEN_3857 = do_replace ? ar_addr : _GEN_3564; // @[playground/src/cache/DCache.scala 259:24 439:26]
  wire [19:0] _GEN_3858 = do_replace ? tag_wdata : _GEN_3565; // @[playground/src/cache/DCache.scala 439:26 183:27]
  wire [63:0] _GEN_3859 = do_replace ? bank_wbdata_0 : _GEN_3566; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3860 = do_replace ? bank_wbdata_1 : _GEN_3567; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3861 = do_replace ? bank_wbdata_2 : _GEN_3568; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3862 = do_replace ? bank_wbdata_3 : _GEN_3569; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3863 = do_replace ? bank_wbdata_4 : _GEN_3570; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3864 = do_replace ? bank_wbdata_5 : _GEN_3571; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3865 = do_replace ? bank_wbdata_6 : _GEN_3572; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3866 = do_replace ? bank_wbdata_7 : _GEN_3573; // @[playground/src/cache/DCache.scala 439:26 166:29]
  wire [63:0] _GEN_3867 = do_replace ? _GEN_295 : _GEN_3574; // @[playground/src/cache/DCache.scala 439:26]
  wire [7:0] _GEN_3868 = do_replace ? _GEN_299 : _GEN_3575; // @[playground/src/cache/DCache.scala 439:26]
  wire [2:0] _GEN_3869 = do_replace ? _GEN_296 : _GEN_3576; // @[playground/src/cache/DCache.scala 439:26]
  wire [7:0] _GEN_3870 = do_replace ? _GEN_298 : _GEN_3579; // @[playground/src/cache/DCache.scala 439:26]
  wire  _GEN_3871 = _T_8 ? _GEN_3583 : _GEN_290; // @[playground/src/cache/DCache.scala 438:29]
  wire  _GEN_3872 = _T_8 ? _GEN_3584 : _GEN_291; // @[playground/src/cache/DCache.scala 438:29]
  wire [2:0] _GEN_3873 = _T_8 ? _GEN_3585 : bank_wbindex; // @[playground/src/cache/DCache.scala 165:29 438:29]
  wire [63:0] _GEN_3874 = _T_8 ? _GEN_3586 : _GEN_297; // @[playground/src/cache/DCache.scala 438:29]
  wire  _GEN_3875 = _T_8 ? _GEN_3587 : _GEN_292; // @[playground/src/cache/DCache.scala 438:29]
  wire  _GEN_3876 = _T_8 ? _GEN_3588 : dirty_0_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3877 = _T_8 ? _GEN_3589 : dirty_0_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3878 = _T_8 ? _GEN_3590 : dirty_1_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3879 = _T_8 ? _GEN_3591 : dirty_1_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3880 = _T_8 ? _GEN_3592 : dirty_2_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3881 = _T_8 ? _GEN_3593 : dirty_2_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3882 = _T_8 ? _GEN_3594 : dirty_3_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3883 = _T_8 ? _GEN_3595 : dirty_3_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3884 = _T_8 ? _GEN_3596 : dirty_4_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3885 = _T_8 ? _GEN_3597 : dirty_4_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3886 = _T_8 ? _GEN_3598 : dirty_5_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3887 = _T_8 ? _GEN_3599 : dirty_5_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3888 = _T_8 ? _GEN_3600 : dirty_6_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3889 = _T_8 ? _GEN_3601 : dirty_6_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3890 = _T_8 ? _GEN_3602 : dirty_7_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3891 = _T_8 ? _GEN_3603 : dirty_7_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3892 = _T_8 ? _GEN_3604 : dirty_8_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3893 = _T_8 ? _GEN_3605 : dirty_8_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3894 = _T_8 ? _GEN_3606 : dirty_9_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3895 = _T_8 ? _GEN_3607 : dirty_9_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3896 = _T_8 ? _GEN_3608 : dirty_10_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3897 = _T_8 ? _GEN_3609 : dirty_10_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3898 = _T_8 ? _GEN_3610 : dirty_11_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3899 = _T_8 ? _GEN_3611 : dirty_11_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3900 = _T_8 ? _GEN_3612 : dirty_12_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3901 = _T_8 ? _GEN_3613 : dirty_12_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3902 = _T_8 ? _GEN_3614 : dirty_13_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3903 = _T_8 ? _GEN_3615 : dirty_13_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3904 = _T_8 ? _GEN_3616 : dirty_14_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3905 = _T_8 ? _GEN_3617 : dirty_14_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3906 = _T_8 ? _GEN_3618 : dirty_15_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3907 = _T_8 ? _GEN_3619 : dirty_15_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3908 = _T_8 ? _GEN_3620 : dirty_16_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3909 = _T_8 ? _GEN_3621 : dirty_16_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3910 = _T_8 ? _GEN_3622 : dirty_17_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3911 = _T_8 ? _GEN_3623 : dirty_17_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3912 = _T_8 ? _GEN_3624 : dirty_18_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3913 = _T_8 ? _GEN_3625 : dirty_18_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3914 = _T_8 ? _GEN_3626 : dirty_19_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3915 = _T_8 ? _GEN_3627 : dirty_19_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3916 = _T_8 ? _GEN_3628 : dirty_20_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3917 = _T_8 ? _GEN_3629 : dirty_20_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3918 = _T_8 ? _GEN_3630 : dirty_21_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3919 = _T_8 ? _GEN_3631 : dirty_21_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3920 = _T_8 ? _GEN_3632 : dirty_22_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3921 = _T_8 ? _GEN_3633 : dirty_22_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3922 = _T_8 ? _GEN_3634 : dirty_23_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3923 = _T_8 ? _GEN_3635 : dirty_23_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3924 = _T_8 ? _GEN_3636 : dirty_24_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3925 = _T_8 ? _GEN_3637 : dirty_24_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3926 = _T_8 ? _GEN_3638 : dirty_25_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3927 = _T_8 ? _GEN_3639 : dirty_25_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3928 = _T_8 ? _GEN_3640 : dirty_26_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3929 = _T_8 ? _GEN_3641 : dirty_26_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3930 = _T_8 ? _GEN_3642 : dirty_27_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3931 = _T_8 ? _GEN_3643 : dirty_27_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3932 = _T_8 ? _GEN_3644 : dirty_28_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3933 = _T_8 ? _GEN_3645 : dirty_28_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3934 = _T_8 ? _GEN_3646 : dirty_29_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3935 = _T_8 ? _GEN_3647 : dirty_29_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3936 = _T_8 ? _GEN_3648 : dirty_30_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3937 = _T_8 ? _GEN_3649 : dirty_30_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3938 = _T_8 ? _GEN_3650 : dirty_31_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3939 = _T_8 ? _GEN_3651 : dirty_31_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3940 = _T_8 ? _GEN_3652 : dirty_32_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3941 = _T_8 ? _GEN_3653 : dirty_32_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3942 = _T_8 ? _GEN_3654 : dirty_33_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3943 = _T_8 ? _GEN_3655 : dirty_33_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3944 = _T_8 ? _GEN_3656 : dirty_34_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3945 = _T_8 ? _GEN_3657 : dirty_34_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3946 = _T_8 ? _GEN_3658 : dirty_35_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3947 = _T_8 ? _GEN_3659 : dirty_35_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3948 = _T_8 ? _GEN_3660 : dirty_36_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3949 = _T_8 ? _GEN_3661 : dirty_36_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3950 = _T_8 ? _GEN_3662 : dirty_37_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3951 = _T_8 ? _GEN_3663 : dirty_37_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3952 = _T_8 ? _GEN_3664 : dirty_38_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3953 = _T_8 ? _GEN_3665 : dirty_38_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3954 = _T_8 ? _GEN_3666 : dirty_39_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3955 = _T_8 ? _GEN_3667 : dirty_39_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3956 = _T_8 ? _GEN_3668 : dirty_40_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3957 = _T_8 ? _GEN_3669 : dirty_40_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3958 = _T_8 ? _GEN_3670 : dirty_41_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3959 = _T_8 ? _GEN_3671 : dirty_41_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3960 = _T_8 ? _GEN_3672 : dirty_42_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3961 = _T_8 ? _GEN_3673 : dirty_42_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3962 = _T_8 ? _GEN_3674 : dirty_43_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3963 = _T_8 ? _GEN_3675 : dirty_43_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3964 = _T_8 ? _GEN_3676 : dirty_44_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3965 = _T_8 ? _GEN_3677 : dirty_44_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3966 = _T_8 ? _GEN_3678 : dirty_45_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3967 = _T_8 ? _GEN_3679 : dirty_45_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3968 = _T_8 ? _GEN_3680 : dirty_46_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3969 = _T_8 ? _GEN_3681 : dirty_46_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3970 = _T_8 ? _GEN_3682 : dirty_47_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3971 = _T_8 ? _GEN_3683 : dirty_47_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3972 = _T_8 ? _GEN_3684 : dirty_48_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3973 = _T_8 ? _GEN_3685 : dirty_48_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3974 = _T_8 ? _GEN_3686 : dirty_49_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3975 = _T_8 ? _GEN_3687 : dirty_49_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3976 = _T_8 ? _GEN_3688 : dirty_50_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3977 = _T_8 ? _GEN_3689 : dirty_50_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3978 = _T_8 ? _GEN_3690 : dirty_51_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3979 = _T_8 ? _GEN_3691 : dirty_51_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3980 = _T_8 ? _GEN_3692 : dirty_52_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3981 = _T_8 ? _GEN_3693 : dirty_52_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3982 = _T_8 ? _GEN_3694 : dirty_53_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3983 = _T_8 ? _GEN_3695 : dirty_53_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3984 = _T_8 ? _GEN_3696 : dirty_54_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3985 = _T_8 ? _GEN_3697 : dirty_54_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3986 = _T_8 ? _GEN_3698 : dirty_55_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3987 = _T_8 ? _GEN_3699 : dirty_55_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3988 = _T_8 ? _GEN_3700 : dirty_56_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3989 = _T_8 ? _GEN_3701 : dirty_56_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3990 = _T_8 ? _GEN_3702 : dirty_57_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3991 = _T_8 ? _GEN_3703 : dirty_57_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3992 = _T_8 ? _GEN_3704 : dirty_58_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3993 = _T_8 ? _GEN_3705 : dirty_58_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3994 = _T_8 ? _GEN_3706 : dirty_59_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3995 = _T_8 ? _GEN_3707 : dirty_59_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3996 = _T_8 ? _GEN_3708 : dirty_60_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3997 = _T_8 ? _GEN_3709 : dirty_60_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3998 = _T_8 ? _GEN_3710 : dirty_61_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_3999 = _T_8 ? _GEN_3711 : dirty_61_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_4000 = _T_8 ? _GEN_3712 : dirty_62_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_4001 = _T_8 ? _GEN_3713 : dirty_62_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_4002 = _T_8 ? _GEN_3714 : dirty_63_0; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_4003 = _T_8 ? _GEN_3715 : dirty_63_1; // @[playground/src/cache/DCache.scala 135:22 438:29]
  wire  _GEN_4004 = _T_8 ? _GEN_3716 : tag_wstrb_0; // @[playground/src/cache/DCache.scala 182:27 438:29]
  wire  _GEN_4005 = _T_8 ? _GEN_3717 : tag_wstrb_1; // @[playground/src/cache/DCache.scala 182:27 438:29]
  wire  _GEN_4006 = _T_8 ? _GEN_3718 : arvalid; // @[playground/src/cache/DCache.scala 260:24 438:29]
  wire  _GEN_4007 = _T_8 ? _GEN_3719 : rready; // @[playground/src/cache/DCache.scala 263:23 438:29]
  wire [7:0] _GEN_4008 = _T_8 ? _GEN_3720 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 160:22 438:29]
  wire [7:0] _GEN_4009 = _T_8 ? _GEN_3721 : burst_wstrb_1; // @[playground/src/cache/DCache.scala 160:22 438:29]
  wire  _GEN_4010 = _T_8 ? _GEN_3722 : valid_0_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4011 = _T_8 ? _GEN_3723 : valid_0_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4012 = _T_8 ? _GEN_3724 : valid_1_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4013 = _T_8 ? _GEN_3725 : valid_1_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4014 = _T_8 ? _GEN_3726 : valid_2_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4015 = _T_8 ? _GEN_3727 : valid_2_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4016 = _T_8 ? _GEN_3728 : valid_3_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4017 = _T_8 ? _GEN_3729 : valid_3_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4018 = _T_8 ? _GEN_3730 : valid_4_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4019 = _T_8 ? _GEN_3731 : valid_4_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4020 = _T_8 ? _GEN_3732 : valid_5_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4021 = _T_8 ? _GEN_3733 : valid_5_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4022 = _T_8 ? _GEN_3734 : valid_6_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4023 = _T_8 ? _GEN_3735 : valid_6_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4024 = _T_8 ? _GEN_3736 : valid_7_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4025 = _T_8 ? _GEN_3737 : valid_7_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4026 = _T_8 ? _GEN_3738 : valid_8_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4027 = _T_8 ? _GEN_3739 : valid_8_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4028 = _T_8 ? _GEN_3740 : valid_9_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4029 = _T_8 ? _GEN_3741 : valid_9_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4030 = _T_8 ? _GEN_3742 : valid_10_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4031 = _T_8 ? _GEN_3743 : valid_10_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4032 = _T_8 ? _GEN_3744 : valid_11_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4033 = _T_8 ? _GEN_3745 : valid_11_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4034 = _T_8 ? _GEN_3746 : valid_12_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4035 = _T_8 ? _GEN_3747 : valid_12_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4036 = _T_8 ? _GEN_3748 : valid_13_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4037 = _T_8 ? _GEN_3749 : valid_13_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4038 = _T_8 ? _GEN_3750 : valid_14_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4039 = _T_8 ? _GEN_3751 : valid_14_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4040 = _T_8 ? _GEN_3752 : valid_15_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4041 = _T_8 ? _GEN_3753 : valid_15_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4042 = _T_8 ? _GEN_3754 : valid_16_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4043 = _T_8 ? _GEN_3755 : valid_16_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4044 = _T_8 ? _GEN_3756 : valid_17_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4045 = _T_8 ? _GEN_3757 : valid_17_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4046 = _T_8 ? _GEN_3758 : valid_18_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4047 = _T_8 ? _GEN_3759 : valid_18_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4048 = _T_8 ? _GEN_3760 : valid_19_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4049 = _T_8 ? _GEN_3761 : valid_19_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4050 = _T_8 ? _GEN_3762 : valid_20_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4051 = _T_8 ? _GEN_3763 : valid_20_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4052 = _T_8 ? _GEN_3764 : valid_21_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4053 = _T_8 ? _GEN_3765 : valid_21_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4054 = _T_8 ? _GEN_3766 : valid_22_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4055 = _T_8 ? _GEN_3767 : valid_22_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4056 = _T_8 ? _GEN_3768 : valid_23_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4057 = _T_8 ? _GEN_3769 : valid_23_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4058 = _T_8 ? _GEN_3770 : valid_24_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4059 = _T_8 ? _GEN_3771 : valid_24_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4060 = _T_8 ? _GEN_3772 : valid_25_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4061 = _T_8 ? _GEN_3773 : valid_25_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4062 = _T_8 ? _GEN_3774 : valid_26_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4063 = _T_8 ? _GEN_3775 : valid_26_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4064 = _T_8 ? _GEN_3776 : valid_27_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4065 = _T_8 ? _GEN_3777 : valid_27_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4066 = _T_8 ? _GEN_3778 : valid_28_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4067 = _T_8 ? _GEN_3779 : valid_28_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4068 = _T_8 ? _GEN_3780 : valid_29_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4069 = _T_8 ? _GEN_3781 : valid_29_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4070 = _T_8 ? _GEN_3782 : valid_30_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4071 = _T_8 ? _GEN_3783 : valid_30_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4072 = _T_8 ? _GEN_3784 : valid_31_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4073 = _T_8 ? _GEN_3785 : valid_31_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4074 = _T_8 ? _GEN_3786 : valid_32_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4075 = _T_8 ? _GEN_3787 : valid_32_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4076 = _T_8 ? _GEN_3788 : valid_33_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4077 = _T_8 ? _GEN_3789 : valid_33_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4078 = _T_8 ? _GEN_3790 : valid_34_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4079 = _T_8 ? _GEN_3791 : valid_34_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4080 = _T_8 ? _GEN_3792 : valid_35_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4081 = _T_8 ? _GEN_3793 : valid_35_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4082 = _T_8 ? _GEN_3794 : valid_36_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4083 = _T_8 ? _GEN_3795 : valid_36_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4084 = _T_8 ? _GEN_3796 : valid_37_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4085 = _T_8 ? _GEN_3797 : valid_37_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4086 = _T_8 ? _GEN_3798 : valid_38_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4087 = _T_8 ? _GEN_3799 : valid_38_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4088 = _T_8 ? _GEN_3800 : valid_39_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4089 = _T_8 ? _GEN_3801 : valid_39_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4090 = _T_8 ? _GEN_3802 : valid_40_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4091 = _T_8 ? _GEN_3803 : valid_40_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4092 = _T_8 ? _GEN_3804 : valid_41_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4093 = _T_8 ? _GEN_3805 : valid_41_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4094 = _T_8 ? _GEN_3806 : valid_42_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4095 = _T_8 ? _GEN_3807 : valid_42_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4096 = _T_8 ? _GEN_3808 : valid_43_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4097 = _T_8 ? _GEN_3809 : valid_43_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4098 = _T_8 ? _GEN_3810 : valid_44_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4099 = _T_8 ? _GEN_3811 : valid_44_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4100 = _T_8 ? _GEN_3812 : valid_45_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4101 = _T_8 ? _GEN_3813 : valid_45_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4102 = _T_8 ? _GEN_3814 : valid_46_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4103 = _T_8 ? _GEN_3815 : valid_46_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4104 = _T_8 ? _GEN_3816 : valid_47_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4105 = _T_8 ? _GEN_3817 : valid_47_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4106 = _T_8 ? _GEN_3818 : valid_48_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4107 = _T_8 ? _GEN_3819 : valid_48_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4108 = _T_8 ? _GEN_3820 : valid_49_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4109 = _T_8 ? _GEN_3821 : valid_49_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4110 = _T_8 ? _GEN_3822 : valid_50_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4111 = _T_8 ? _GEN_3823 : valid_50_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4112 = _T_8 ? _GEN_3824 : valid_51_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4113 = _T_8 ? _GEN_3825 : valid_51_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4114 = _T_8 ? _GEN_3826 : valid_52_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4115 = _T_8 ? _GEN_3827 : valid_52_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4116 = _T_8 ? _GEN_3828 : valid_53_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4117 = _T_8 ? _GEN_3829 : valid_53_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4118 = _T_8 ? _GEN_3830 : valid_54_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4119 = _T_8 ? _GEN_3831 : valid_54_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4120 = _T_8 ? _GEN_3832 : valid_55_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4121 = _T_8 ? _GEN_3833 : valid_55_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4122 = _T_8 ? _GEN_3834 : valid_56_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4123 = _T_8 ? _GEN_3835 : valid_56_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4124 = _T_8 ? _GEN_3836 : valid_57_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4125 = _T_8 ? _GEN_3837 : valid_57_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4126 = _T_8 ? _GEN_3838 : valid_58_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4127 = _T_8 ? _GEN_3839 : valid_58_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4128 = _T_8 ? _GEN_3840 : valid_59_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4129 = _T_8 ? _GEN_3841 : valid_59_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4130 = _T_8 ? _GEN_3842 : valid_60_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4131 = _T_8 ? _GEN_3843 : valid_60_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4132 = _T_8 ? _GEN_3844 : valid_61_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4133 = _T_8 ? _GEN_3845 : valid_61_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4134 = _T_8 ? _GEN_3846 : valid_62_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4135 = _T_8 ? _GEN_3847 : valid_62_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4136 = _T_8 ? _GEN_3848 : valid_63_0; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4137 = _T_8 ? _GEN_3849 : valid_63_1; // @[playground/src/cache/DCache.scala 134:22 438:29]
  wire  _GEN_4138 = _T_8 ? _GEN_3850 : do_replace; // @[playground/src/cache/DCache.scala 438:29 170:30]
  wire  _GEN_4139 = _T_8 ? _GEN_3851 : ptw_scratch_replace; // @[playground/src/cache/DCache.scala 101:28 438:29]
  wire [2:0] _GEN_4140 = _T_8 ? _GEN_3852 : state; // @[playground/src/cache/DCache.scala 438:29 90:94]
  wire  _GEN_4141 = _T_8 ? _GEN_3853 : ptw_scratch_dcache_wait; // @[playground/src/cache/DCache.scala 101:28 438:29]
  wire  _GEN_4142 = _T_8 ? _GEN_3854 : readsram; // @[playground/src/cache/DCache.scala 148:25 438:29]
  wire [7:0] _GEN_4143 = _T_8 ? _GEN_3855 : ar_len; // @[playground/src/cache/DCache.scala 259:24 438:29]
  wire [2:0] _GEN_4144 = _T_8 ? _GEN_3856 : ar_size; // @[playground/src/cache/DCache.scala 259:24 438:29]
  wire [31:0] _GEN_4145 = _T_8 ? _GEN_3857 : ar_addr; // @[playground/src/cache/DCache.scala 259:24 438:29]
  wire [19:0] _GEN_4146 = _T_8 ? _GEN_3858 : tag_wdata; // @[playground/src/cache/DCache.scala 183:27 438:29]
  wire [63:0] _GEN_4147 = _T_8 ? _GEN_3859 : bank_wbdata_0; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4148 = _T_8 ? _GEN_3860 : bank_wbdata_1; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4149 = _T_8 ? _GEN_3861 : bank_wbdata_2; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4150 = _T_8 ? _GEN_3862 : bank_wbdata_3; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4151 = _T_8 ? _GEN_3863 : bank_wbdata_4; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4152 = _T_8 ? _GEN_3864 : bank_wbdata_5; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4153 = _T_8 ? _GEN_3865 : bank_wbdata_6; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4154 = _T_8 ? _GEN_3866 : bank_wbdata_7; // @[playground/src/cache/DCache.scala 166:29 438:29]
  wire [63:0] _GEN_4155 = _T_8 ? _GEN_3867 : _GEN_295; // @[playground/src/cache/DCache.scala 438:29]
  wire [7:0] _GEN_4156 = _T_8 ? _GEN_3868 : _GEN_299; // @[playground/src/cache/DCache.scala 438:29]
  wire [2:0] _GEN_4157 = _T_8 ? _GEN_3869 : _GEN_296; // @[playground/src/cache/DCache.scala 438:29]
  wire [7:0] _GEN_4158 = _T_8 ? _GEN_3870 : _GEN_298; // @[playground/src/cache/DCache.scala 438:29]
  wire  _GEN_4159 = io_cpu_complete_single_request ? 1'h0 : 1'h1; // @[playground/src/cache/DCache.scala 534:32 535:44 536:33]
  wire  _GEN_4160 = io_cpu_complete_single_request ? 1'h0 : access_fault; // @[playground/src/cache/DCache.scala 277:29 535:44 537:33]
  wire  _GEN_4161 = io_cpu_complete_single_request ? 1'h0 : page_fault; // @[playground/src/cache/DCache.scala 278:29 535:44 538:33]
  wire [2:0] _GEN_4162 = io_cpu_complete_single_request ? 3'h0 : state; // @[playground/src/cache/DCache.scala 535:44 539:33 90:94]
  wire [2:0] _GEN_4163 = io_cpu_tlb_hit ? 3'h0 : state; // @[playground/src/cache/DCache.scala 551:30 552:17 90:94]
  wire  _GEN_4164 = io_cpu_tlb_page_fault | page_fault; // @[playground/src/cache/DCache.scala 547:41 548:20 278:29]
  wire [2:0] _GEN_4165 = io_cpu_tlb_page_fault ? 3'h4 : _GEN_4163; // @[playground/src/cache/DCache.scala 547:41 549:20]
  wire  _GEN_4169 = 3'h5 == state & _io_cpu_tlb_ptw_vpn_ready_T; // @[playground/src/cache/DCache.scala 316:17 107:28 543:32]
  wire [2:0] _GEN_4171 = 3'h5 == state ? _GEN_4165 : state; // @[playground/src/cache/DCache.scala 316:17 90:94]
  wire  _GEN_4172 = 3'h5 == state ? _GEN_4164 : page_fault; // @[playground/src/cache/DCache.scala 316:17 278:29]
  wire  _GEN_4173 = 3'h4 == state ? _io_cpu_tlb_ptw_vpn_ready_T : _GEN_4169; // @[playground/src/cache/DCache.scala 316:17 533:32]
  wire  _GEN_4174 = 3'h4 == state ? _GEN_4159 : ptw_scratch_dcache_wait; // @[playground/src/cache/DCache.scala 316:17 101:28]
  wire  _GEN_4175 = 3'h4 == state ? _GEN_4160 : access_fault; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4176 = 3'h4 == state ? _GEN_4161 : _GEN_4172; // @[playground/src/cache/DCache.scala 316:17]
  wire [2:0] _GEN_4177 = 3'h4 == state ? _GEN_4162 : _GEN_4171; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4178 = 3'h3 == state ? _GEN_3871 : _GEN_290; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4179 = 3'h3 == state ? _GEN_3872 : _GEN_291; // @[playground/src/cache/DCache.scala 316:17]
  wire [2:0] _GEN_4180 = 3'h3 == state ? _GEN_3873 : bank_wbindex; // @[playground/src/cache/DCache.scala 316:17 165:29]
  wire [63:0] _GEN_4181 = 3'h3 == state ? _GEN_3874 : _GEN_297; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4182 = 3'h3 == state ? _GEN_3875 : _GEN_292; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4183 = 3'h3 == state ? _GEN_3876 : dirty_0_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4184 = 3'h3 == state ? _GEN_3877 : dirty_0_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4185 = 3'h3 == state ? _GEN_3878 : dirty_1_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4186 = 3'h3 == state ? _GEN_3879 : dirty_1_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4187 = 3'h3 == state ? _GEN_3880 : dirty_2_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4188 = 3'h3 == state ? _GEN_3881 : dirty_2_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4189 = 3'h3 == state ? _GEN_3882 : dirty_3_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4190 = 3'h3 == state ? _GEN_3883 : dirty_3_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4191 = 3'h3 == state ? _GEN_3884 : dirty_4_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4192 = 3'h3 == state ? _GEN_3885 : dirty_4_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4193 = 3'h3 == state ? _GEN_3886 : dirty_5_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4194 = 3'h3 == state ? _GEN_3887 : dirty_5_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4195 = 3'h3 == state ? _GEN_3888 : dirty_6_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4196 = 3'h3 == state ? _GEN_3889 : dirty_6_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4197 = 3'h3 == state ? _GEN_3890 : dirty_7_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4198 = 3'h3 == state ? _GEN_3891 : dirty_7_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4199 = 3'h3 == state ? _GEN_3892 : dirty_8_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4200 = 3'h3 == state ? _GEN_3893 : dirty_8_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4201 = 3'h3 == state ? _GEN_3894 : dirty_9_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4202 = 3'h3 == state ? _GEN_3895 : dirty_9_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4203 = 3'h3 == state ? _GEN_3896 : dirty_10_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4204 = 3'h3 == state ? _GEN_3897 : dirty_10_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4205 = 3'h3 == state ? _GEN_3898 : dirty_11_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4206 = 3'h3 == state ? _GEN_3899 : dirty_11_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4207 = 3'h3 == state ? _GEN_3900 : dirty_12_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4208 = 3'h3 == state ? _GEN_3901 : dirty_12_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4209 = 3'h3 == state ? _GEN_3902 : dirty_13_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4210 = 3'h3 == state ? _GEN_3903 : dirty_13_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4211 = 3'h3 == state ? _GEN_3904 : dirty_14_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4212 = 3'h3 == state ? _GEN_3905 : dirty_14_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4213 = 3'h3 == state ? _GEN_3906 : dirty_15_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4214 = 3'h3 == state ? _GEN_3907 : dirty_15_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4215 = 3'h3 == state ? _GEN_3908 : dirty_16_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4216 = 3'h3 == state ? _GEN_3909 : dirty_16_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4217 = 3'h3 == state ? _GEN_3910 : dirty_17_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4218 = 3'h3 == state ? _GEN_3911 : dirty_17_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4219 = 3'h3 == state ? _GEN_3912 : dirty_18_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4220 = 3'h3 == state ? _GEN_3913 : dirty_18_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4221 = 3'h3 == state ? _GEN_3914 : dirty_19_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4222 = 3'h3 == state ? _GEN_3915 : dirty_19_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4223 = 3'h3 == state ? _GEN_3916 : dirty_20_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4224 = 3'h3 == state ? _GEN_3917 : dirty_20_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4225 = 3'h3 == state ? _GEN_3918 : dirty_21_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4226 = 3'h3 == state ? _GEN_3919 : dirty_21_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4227 = 3'h3 == state ? _GEN_3920 : dirty_22_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4228 = 3'h3 == state ? _GEN_3921 : dirty_22_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4229 = 3'h3 == state ? _GEN_3922 : dirty_23_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4230 = 3'h3 == state ? _GEN_3923 : dirty_23_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4231 = 3'h3 == state ? _GEN_3924 : dirty_24_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4232 = 3'h3 == state ? _GEN_3925 : dirty_24_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4233 = 3'h3 == state ? _GEN_3926 : dirty_25_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4234 = 3'h3 == state ? _GEN_3927 : dirty_25_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4235 = 3'h3 == state ? _GEN_3928 : dirty_26_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4236 = 3'h3 == state ? _GEN_3929 : dirty_26_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4237 = 3'h3 == state ? _GEN_3930 : dirty_27_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4238 = 3'h3 == state ? _GEN_3931 : dirty_27_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4239 = 3'h3 == state ? _GEN_3932 : dirty_28_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4240 = 3'h3 == state ? _GEN_3933 : dirty_28_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4241 = 3'h3 == state ? _GEN_3934 : dirty_29_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4242 = 3'h3 == state ? _GEN_3935 : dirty_29_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4243 = 3'h3 == state ? _GEN_3936 : dirty_30_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4244 = 3'h3 == state ? _GEN_3937 : dirty_30_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4245 = 3'h3 == state ? _GEN_3938 : dirty_31_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4246 = 3'h3 == state ? _GEN_3939 : dirty_31_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4247 = 3'h3 == state ? _GEN_3940 : dirty_32_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4248 = 3'h3 == state ? _GEN_3941 : dirty_32_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4249 = 3'h3 == state ? _GEN_3942 : dirty_33_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4250 = 3'h3 == state ? _GEN_3943 : dirty_33_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4251 = 3'h3 == state ? _GEN_3944 : dirty_34_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4252 = 3'h3 == state ? _GEN_3945 : dirty_34_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4253 = 3'h3 == state ? _GEN_3946 : dirty_35_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4254 = 3'h3 == state ? _GEN_3947 : dirty_35_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4255 = 3'h3 == state ? _GEN_3948 : dirty_36_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4256 = 3'h3 == state ? _GEN_3949 : dirty_36_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4257 = 3'h3 == state ? _GEN_3950 : dirty_37_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4258 = 3'h3 == state ? _GEN_3951 : dirty_37_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4259 = 3'h3 == state ? _GEN_3952 : dirty_38_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4260 = 3'h3 == state ? _GEN_3953 : dirty_38_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4261 = 3'h3 == state ? _GEN_3954 : dirty_39_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4262 = 3'h3 == state ? _GEN_3955 : dirty_39_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4263 = 3'h3 == state ? _GEN_3956 : dirty_40_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4264 = 3'h3 == state ? _GEN_3957 : dirty_40_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4265 = 3'h3 == state ? _GEN_3958 : dirty_41_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4266 = 3'h3 == state ? _GEN_3959 : dirty_41_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4267 = 3'h3 == state ? _GEN_3960 : dirty_42_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4268 = 3'h3 == state ? _GEN_3961 : dirty_42_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4269 = 3'h3 == state ? _GEN_3962 : dirty_43_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4270 = 3'h3 == state ? _GEN_3963 : dirty_43_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4271 = 3'h3 == state ? _GEN_3964 : dirty_44_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4272 = 3'h3 == state ? _GEN_3965 : dirty_44_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4273 = 3'h3 == state ? _GEN_3966 : dirty_45_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4274 = 3'h3 == state ? _GEN_3967 : dirty_45_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4275 = 3'h3 == state ? _GEN_3968 : dirty_46_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4276 = 3'h3 == state ? _GEN_3969 : dirty_46_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4277 = 3'h3 == state ? _GEN_3970 : dirty_47_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4278 = 3'h3 == state ? _GEN_3971 : dirty_47_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4279 = 3'h3 == state ? _GEN_3972 : dirty_48_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4280 = 3'h3 == state ? _GEN_3973 : dirty_48_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4281 = 3'h3 == state ? _GEN_3974 : dirty_49_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4282 = 3'h3 == state ? _GEN_3975 : dirty_49_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4283 = 3'h3 == state ? _GEN_3976 : dirty_50_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4284 = 3'h3 == state ? _GEN_3977 : dirty_50_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4285 = 3'h3 == state ? _GEN_3978 : dirty_51_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4286 = 3'h3 == state ? _GEN_3979 : dirty_51_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4287 = 3'h3 == state ? _GEN_3980 : dirty_52_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4288 = 3'h3 == state ? _GEN_3981 : dirty_52_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4289 = 3'h3 == state ? _GEN_3982 : dirty_53_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4290 = 3'h3 == state ? _GEN_3983 : dirty_53_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4291 = 3'h3 == state ? _GEN_3984 : dirty_54_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4292 = 3'h3 == state ? _GEN_3985 : dirty_54_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4293 = 3'h3 == state ? _GEN_3986 : dirty_55_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4294 = 3'h3 == state ? _GEN_3987 : dirty_55_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4295 = 3'h3 == state ? _GEN_3988 : dirty_56_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4296 = 3'h3 == state ? _GEN_3989 : dirty_56_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4297 = 3'h3 == state ? _GEN_3990 : dirty_57_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4298 = 3'h3 == state ? _GEN_3991 : dirty_57_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4299 = 3'h3 == state ? _GEN_3992 : dirty_58_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4300 = 3'h3 == state ? _GEN_3993 : dirty_58_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4301 = 3'h3 == state ? _GEN_3994 : dirty_59_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4302 = 3'h3 == state ? _GEN_3995 : dirty_59_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4303 = 3'h3 == state ? _GEN_3996 : dirty_60_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4304 = 3'h3 == state ? _GEN_3997 : dirty_60_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4305 = 3'h3 == state ? _GEN_3998 : dirty_61_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4306 = 3'h3 == state ? _GEN_3999 : dirty_61_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4307 = 3'h3 == state ? _GEN_4000 : dirty_62_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4308 = 3'h3 == state ? _GEN_4001 : dirty_62_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4309 = 3'h3 == state ? _GEN_4002 : dirty_63_0; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4310 = 3'h3 == state ? _GEN_4003 : dirty_63_1; // @[playground/src/cache/DCache.scala 316:17 135:22]
  wire  _GEN_4311 = 3'h3 == state ? _GEN_4004 : tag_wstrb_0; // @[playground/src/cache/DCache.scala 316:17 182:27]
  wire  _GEN_4312 = 3'h3 == state ? _GEN_4005 : tag_wstrb_1; // @[playground/src/cache/DCache.scala 316:17 182:27]
  wire  _GEN_4313 = 3'h3 == state ? _GEN_4006 : arvalid; // @[playground/src/cache/DCache.scala 316:17 260:24]
  wire  _GEN_4314 = 3'h3 == state ? _GEN_4007 : rready; // @[playground/src/cache/DCache.scala 316:17 263:23]
  wire [7:0] _GEN_4315 = 3'h3 == state ? _GEN_4008 : burst_wstrb_0; // @[playground/src/cache/DCache.scala 316:17 160:22]
  wire [7:0] _GEN_4316 = 3'h3 == state ? _GEN_4009 : burst_wstrb_1; // @[playground/src/cache/DCache.scala 316:17 160:22]
  wire  _GEN_4317 = 3'h3 == state ? _GEN_4010 : valid_0_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4318 = 3'h3 == state ? _GEN_4011 : valid_0_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4319 = 3'h3 == state ? _GEN_4012 : valid_1_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4320 = 3'h3 == state ? _GEN_4013 : valid_1_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4321 = 3'h3 == state ? _GEN_4014 : valid_2_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4322 = 3'h3 == state ? _GEN_4015 : valid_2_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4323 = 3'h3 == state ? _GEN_4016 : valid_3_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4324 = 3'h3 == state ? _GEN_4017 : valid_3_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4325 = 3'h3 == state ? _GEN_4018 : valid_4_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4326 = 3'h3 == state ? _GEN_4019 : valid_4_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4327 = 3'h3 == state ? _GEN_4020 : valid_5_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4328 = 3'h3 == state ? _GEN_4021 : valid_5_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4329 = 3'h3 == state ? _GEN_4022 : valid_6_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4330 = 3'h3 == state ? _GEN_4023 : valid_6_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4331 = 3'h3 == state ? _GEN_4024 : valid_7_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4332 = 3'h3 == state ? _GEN_4025 : valid_7_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4333 = 3'h3 == state ? _GEN_4026 : valid_8_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4334 = 3'h3 == state ? _GEN_4027 : valid_8_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4335 = 3'h3 == state ? _GEN_4028 : valid_9_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4336 = 3'h3 == state ? _GEN_4029 : valid_9_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4337 = 3'h3 == state ? _GEN_4030 : valid_10_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4338 = 3'h3 == state ? _GEN_4031 : valid_10_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4339 = 3'h3 == state ? _GEN_4032 : valid_11_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4340 = 3'h3 == state ? _GEN_4033 : valid_11_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4341 = 3'h3 == state ? _GEN_4034 : valid_12_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4342 = 3'h3 == state ? _GEN_4035 : valid_12_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4343 = 3'h3 == state ? _GEN_4036 : valid_13_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4344 = 3'h3 == state ? _GEN_4037 : valid_13_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4345 = 3'h3 == state ? _GEN_4038 : valid_14_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4346 = 3'h3 == state ? _GEN_4039 : valid_14_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4347 = 3'h3 == state ? _GEN_4040 : valid_15_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4348 = 3'h3 == state ? _GEN_4041 : valid_15_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4349 = 3'h3 == state ? _GEN_4042 : valid_16_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4350 = 3'h3 == state ? _GEN_4043 : valid_16_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4351 = 3'h3 == state ? _GEN_4044 : valid_17_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4352 = 3'h3 == state ? _GEN_4045 : valid_17_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4353 = 3'h3 == state ? _GEN_4046 : valid_18_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4354 = 3'h3 == state ? _GEN_4047 : valid_18_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4355 = 3'h3 == state ? _GEN_4048 : valid_19_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4356 = 3'h3 == state ? _GEN_4049 : valid_19_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4357 = 3'h3 == state ? _GEN_4050 : valid_20_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4358 = 3'h3 == state ? _GEN_4051 : valid_20_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4359 = 3'h3 == state ? _GEN_4052 : valid_21_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4360 = 3'h3 == state ? _GEN_4053 : valid_21_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4361 = 3'h3 == state ? _GEN_4054 : valid_22_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4362 = 3'h3 == state ? _GEN_4055 : valid_22_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4363 = 3'h3 == state ? _GEN_4056 : valid_23_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4364 = 3'h3 == state ? _GEN_4057 : valid_23_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4365 = 3'h3 == state ? _GEN_4058 : valid_24_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4366 = 3'h3 == state ? _GEN_4059 : valid_24_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4367 = 3'h3 == state ? _GEN_4060 : valid_25_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4368 = 3'h3 == state ? _GEN_4061 : valid_25_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4369 = 3'h3 == state ? _GEN_4062 : valid_26_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4370 = 3'h3 == state ? _GEN_4063 : valid_26_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4371 = 3'h3 == state ? _GEN_4064 : valid_27_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4372 = 3'h3 == state ? _GEN_4065 : valid_27_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4373 = 3'h3 == state ? _GEN_4066 : valid_28_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4374 = 3'h3 == state ? _GEN_4067 : valid_28_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4375 = 3'h3 == state ? _GEN_4068 : valid_29_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4376 = 3'h3 == state ? _GEN_4069 : valid_29_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4377 = 3'h3 == state ? _GEN_4070 : valid_30_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4378 = 3'h3 == state ? _GEN_4071 : valid_30_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4379 = 3'h3 == state ? _GEN_4072 : valid_31_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4380 = 3'h3 == state ? _GEN_4073 : valid_31_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4381 = 3'h3 == state ? _GEN_4074 : valid_32_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4382 = 3'h3 == state ? _GEN_4075 : valid_32_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4383 = 3'h3 == state ? _GEN_4076 : valid_33_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4384 = 3'h3 == state ? _GEN_4077 : valid_33_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4385 = 3'h3 == state ? _GEN_4078 : valid_34_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4386 = 3'h3 == state ? _GEN_4079 : valid_34_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4387 = 3'h3 == state ? _GEN_4080 : valid_35_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4388 = 3'h3 == state ? _GEN_4081 : valid_35_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4389 = 3'h3 == state ? _GEN_4082 : valid_36_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4390 = 3'h3 == state ? _GEN_4083 : valid_36_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4391 = 3'h3 == state ? _GEN_4084 : valid_37_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4392 = 3'h3 == state ? _GEN_4085 : valid_37_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4393 = 3'h3 == state ? _GEN_4086 : valid_38_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4394 = 3'h3 == state ? _GEN_4087 : valid_38_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4395 = 3'h3 == state ? _GEN_4088 : valid_39_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4396 = 3'h3 == state ? _GEN_4089 : valid_39_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4397 = 3'h3 == state ? _GEN_4090 : valid_40_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4398 = 3'h3 == state ? _GEN_4091 : valid_40_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4399 = 3'h3 == state ? _GEN_4092 : valid_41_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4400 = 3'h3 == state ? _GEN_4093 : valid_41_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4401 = 3'h3 == state ? _GEN_4094 : valid_42_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4402 = 3'h3 == state ? _GEN_4095 : valid_42_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4403 = 3'h3 == state ? _GEN_4096 : valid_43_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4404 = 3'h3 == state ? _GEN_4097 : valid_43_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4405 = 3'h3 == state ? _GEN_4098 : valid_44_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4406 = 3'h3 == state ? _GEN_4099 : valid_44_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4407 = 3'h3 == state ? _GEN_4100 : valid_45_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4408 = 3'h3 == state ? _GEN_4101 : valid_45_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4409 = 3'h3 == state ? _GEN_4102 : valid_46_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4410 = 3'h3 == state ? _GEN_4103 : valid_46_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4411 = 3'h3 == state ? _GEN_4104 : valid_47_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4412 = 3'h3 == state ? _GEN_4105 : valid_47_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4413 = 3'h3 == state ? _GEN_4106 : valid_48_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4414 = 3'h3 == state ? _GEN_4107 : valid_48_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4415 = 3'h3 == state ? _GEN_4108 : valid_49_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4416 = 3'h3 == state ? _GEN_4109 : valid_49_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4417 = 3'h3 == state ? _GEN_4110 : valid_50_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4418 = 3'h3 == state ? _GEN_4111 : valid_50_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4419 = 3'h3 == state ? _GEN_4112 : valid_51_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4420 = 3'h3 == state ? _GEN_4113 : valid_51_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4421 = 3'h3 == state ? _GEN_4114 : valid_52_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4422 = 3'h3 == state ? _GEN_4115 : valid_52_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4423 = 3'h3 == state ? _GEN_4116 : valid_53_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4424 = 3'h3 == state ? _GEN_4117 : valid_53_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4425 = 3'h3 == state ? _GEN_4118 : valid_54_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4426 = 3'h3 == state ? _GEN_4119 : valid_54_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4427 = 3'h3 == state ? _GEN_4120 : valid_55_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4428 = 3'h3 == state ? _GEN_4121 : valid_55_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4429 = 3'h3 == state ? _GEN_4122 : valid_56_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4430 = 3'h3 == state ? _GEN_4123 : valid_56_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4431 = 3'h3 == state ? _GEN_4124 : valid_57_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4432 = 3'h3 == state ? _GEN_4125 : valid_57_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4433 = 3'h3 == state ? _GEN_4126 : valid_58_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4434 = 3'h3 == state ? _GEN_4127 : valid_58_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4435 = 3'h3 == state ? _GEN_4128 : valid_59_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4436 = 3'h3 == state ? _GEN_4129 : valid_59_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4437 = 3'h3 == state ? _GEN_4130 : valid_60_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4438 = 3'h3 == state ? _GEN_4131 : valid_60_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4439 = 3'h3 == state ? _GEN_4132 : valid_61_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4440 = 3'h3 == state ? _GEN_4133 : valid_61_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4441 = 3'h3 == state ? _GEN_4134 : valid_62_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4442 = 3'h3 == state ? _GEN_4135 : valid_62_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4443 = 3'h3 == state ? _GEN_4136 : valid_63_0; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4444 = 3'h3 == state ? _GEN_4137 : valid_63_1; // @[playground/src/cache/DCache.scala 316:17 134:22]
  wire  _GEN_4445 = 3'h3 == state ? _GEN_4138 : do_replace; // @[playground/src/cache/DCache.scala 316:17 170:30]
  wire  _GEN_4446 = 3'h3 == state ? _GEN_4139 : ptw_scratch_replace; // @[playground/src/cache/DCache.scala 316:17 101:28]
  wire [2:0] _GEN_4447 = 3'h3 == state ? _GEN_4140 : _GEN_4177; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4448 = 3'h3 == state ? _GEN_4141 : _GEN_4174; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4449 = 3'h3 == state ? _GEN_4142 : readsram; // @[playground/src/cache/DCache.scala 316:17 148:25]
  wire [7:0] _GEN_4450 = 3'h3 == state ? _GEN_4143 : ar_len; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [2:0] _GEN_4451 = 3'h3 == state ? _GEN_4144 : ar_size; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [31:0] _GEN_4452 = 3'h3 == state ? _GEN_4145 : ar_addr; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [19:0] _GEN_4453 = 3'h3 == state ? _GEN_4146 : tag_wdata; // @[playground/src/cache/DCache.scala 316:17 183:27]
  wire [63:0] _GEN_4454 = 3'h3 == state ? _GEN_4147 : bank_wbdata_0; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4455 = 3'h3 == state ? _GEN_4148 : bank_wbdata_1; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4456 = 3'h3 == state ? _GEN_4149 : bank_wbdata_2; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4457 = 3'h3 == state ? _GEN_4150 : bank_wbdata_3; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4458 = 3'h3 == state ? _GEN_4151 : bank_wbdata_4; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4459 = 3'h3 == state ? _GEN_4152 : bank_wbdata_5; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4460 = 3'h3 == state ? _GEN_4153 : bank_wbdata_6; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4461 = 3'h3 == state ? _GEN_4154 : bank_wbdata_7; // @[playground/src/cache/DCache.scala 316:17 166:29]
  wire [63:0] _GEN_4462 = 3'h3 == state ? _GEN_4155 : _GEN_295; // @[playground/src/cache/DCache.scala 316:17]
  wire [7:0] _GEN_4463 = 3'h3 == state ? _GEN_4156 : _GEN_299; // @[playground/src/cache/DCache.scala 316:17]
  wire [2:0] _GEN_4464 = 3'h3 == state ? _GEN_4157 : _GEN_296; // @[playground/src/cache/DCache.scala 316:17]
  wire [7:0] _GEN_4465 = 3'h3 == state ? _GEN_4158 : _GEN_298; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4466 = 3'h3 == state ? 1'h0 : _GEN_4173; // @[playground/src/cache/DCache.scala 316:17 107:28]
  wire  _GEN_4467 = 3'h3 == state ? access_fault : _GEN_4175; // @[playground/src/cache/DCache.scala 316:17 277:29]
  wire  _GEN_4468 = 3'h3 == state ? page_fault : _GEN_4176; // @[playground/src/cache/DCache.scala 316:17 278:29]
  wire [63:0] _GEN_4604 = 3'h2 == state ? _GEN_2372 : _GEN_4462; // @[playground/src/cache/DCache.scala 316:17]
  wire [2:0] _GEN_4608 = 3'h2 == state ? _GEN_2376 : _GEN_4447; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4611 = 3'h2 == state ? arvalid : _GEN_4313; // @[playground/src/cache/DCache.scala 316:17 260:24]
  wire  _GEN_4612 = 3'h2 == state ? rready : _GEN_4314; // @[playground/src/cache/DCache.scala 316:17 263:23]
  wire  _GEN_4744 = 3'h2 == state ? ptw_scratch_replace : _GEN_4446; // @[playground/src/cache/DCache.scala 316:17 101:28]
  wire [7:0] _GEN_4746 = 3'h2 == state ? ar_len : _GEN_4450; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [2:0] _GEN_4747 = 3'h2 == state ? ar_size : _GEN_4451; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [31:0] _GEN_4748 = 3'h2 == state ? ar_addr : _GEN_4452; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire  _GEN_4758 = 3'h2 == state ? 1'h0 : _GEN_4466; // @[playground/src/cache/DCache.scala 316:17 107:28]
  wire  _GEN_4761 = 3'h1 == state ? _GEN_1860 : _GEN_4611; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_4762 = 3'h1 == state ? _GEN_1861 : _GEN_4612; // @[playground/src/cache/DCache.scala 316:17]
  wire [2:0] _GEN_4765 = 3'h1 == state ? _GEN_1864 : _GEN_4608; // @[playground/src/cache/DCache.scala 316:17]
  wire [63:0] _GEN_4901 = 3'h1 == state ? _GEN_295 : _GEN_4604; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_5038 = 3'h1 == state ? ptw_scratch_replace : _GEN_4744; // @[playground/src/cache/DCache.scala 316:17 101:28]
  wire [7:0] _GEN_5040 = 3'h1 == state ? ar_len : _GEN_4746; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [2:0] _GEN_5041 = 3'h1 == state ? ar_size : _GEN_4747; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire [31:0] _GEN_5042 = 3'h1 == state ? ar_addr : _GEN_4748; // @[playground/src/cache/DCache.scala 316:17 259:24]
  wire  _GEN_5052 = 3'h1 == state ? 1'h0 : _GEN_4758; // @[playground/src/cache/DCache.scala 316:17 107:28]
  wire [2:0] _GEN_5056 = 3'h0 == state ? _GEN_1654 : _GEN_4765; // @[playground/src/cache/DCache.scala 316:17]
  wire [7:0] _GEN_5059 = 3'h0 == state ? _GEN_1657 : 8'h0; // @[playground/src/cache/DCache.scala 316:17 156:26]
  wire [31:0] _GEN_5062 = 3'h0 == state ? _GEN_1660 : _GEN_5042; // @[playground/src/cache/DCache.scala 316:17]
  wire [7:0] _GEN_5063 = 3'h0 == state ? _GEN_1661 : _GEN_5040; // @[playground/src/cache/DCache.scala 316:17]
  wire [7:0] _GEN_5064 = 3'h0 == state ? _GEN_1662 : {{5'd0}, _GEN_5041}; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_5065 = 3'h0 == state ? _GEN_1663 : _GEN_4761; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_5066 = 3'h0 == state ? _GEN_1664 : _GEN_4762; // @[playground/src/cache/DCache.scala 316:17]
  wire [63:0] _GEN_5268 = 3'h0 == state ? _GEN_295 : _GEN_4901; // @[playground/src/cache/DCache.scala 316:17]
  wire  _GEN_5405 = 3'h0 == state ? ptw_scratch_replace : _GEN_5038; // @[playground/src/cache/DCache.scala 316:17 101:28]
  wire [19:0] satp_ppn = io_cpu_tlb_csr_satp[19:0]; // @[playground/src/cache/DCache.scala 560:49]
  wire  mstatus_sum = io_cpu_tlb_csr_mstatus[18]; // @[playground/src/cache/DCache.scala 561:52]
  wire  mstatus_mxr = io_cpu_tlb_csr_mstatus[19]; // @[playground/src/cache/DCache.scala 561:52]
  wire [1:0] mode = io_cpu_tlb_access_type == 2'h0 ? io_cpu_tlb_csr_imode : io_cpu_tlb_csr_dmode; // @[playground/src/cache/DCache.scala 562:24]
  reg [19:0] pte_ppn; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_d; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_a; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_g; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_u; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_x; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_w; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_r; // @[playground/src/cache/DCache.scala 569:28]
  reg  pte_flag_v; // @[playground/src/cache/DCache.scala 569:28]
  wire  _T_50 = io_cpu_tlb_ptw_vpn_ready & io_cpu_tlb_ptw_vpn_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _GEN_5419 = pte_uncached | _GEN_5065; // @[playground/src/cache/DCache.scala 622:26 623:19]
  wire [7:0] _GEN_5421 = pte_uncached ? 8'h3 : _GEN_5064; // @[playground/src/cache/DCache.scala 622:26 625:19]
  wire  _GEN_5423 = pte_uncached | _GEN_5066; // @[playground/src/cache/DCache.scala 622:26 627:19]
  wire [5:0] _GEN_5425 = pte_uncached ? _bank_raddr_T_2 : ptw_addr_index; // @[playground/src/cache/DCache.scala 218:14 622:26 630:31]
  wire  _GEN_5431 = pte_uncached & _GEN_5405; // @[playground/src/cache/DCache.scala 622:26 635:31]
  wire [63:0] _GEN_5561 = 3'h0 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_0_1 : data_0_0; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5562 = 3'h1 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_1_0 : _GEN_5561; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5563 = 3'h1 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_1_1 : _GEN_5562; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5564 = 3'h2 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_2_0 : _GEN_5563; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5565 = 3'h2 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_2_1 : _GEN_5564; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5566 = 3'h3 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_3_0 : _GEN_5565; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5567 = 3'h3 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_3_1 : _GEN_5566; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5568 = 3'h4 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_4_0 : _GEN_5567; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5569 = 3'h4 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_4_1 : _GEN_5568; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5570 = 3'h5 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_5_0 : _GEN_5569; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5571 = 3'h5 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_5_1 : _GEN_5570; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5572 = 3'h6 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_6_0 : _GEN_5571; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5573 = 3'h6 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_6_1 : _GEN_5572; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5574 = 3'h7 == ptw_scratch_paddr_offset[5:3] & _GEN_5964 ? data_7_0 : _GEN_5573; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire [63:0] _GEN_5575 = 3'h7 == ptw_scratch_paddr_offset[5:3] & tag_compare_valid_1 ? data_7_1 : _GEN_5574; // @[playground/src/cache/DCache.scala 649:{102,102}]
  wire  pte_temp_flag_v = _GEN_5575[0]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_r = _GEN_5575[1]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_w = _GEN_5575[2]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_x = _GEN_5575[3]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_u = _GEN_5575[4]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_g = _GEN_5575[5]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_a = _GEN_5575[6]; // @[playground/src/cache/DCache.scala 649:102]
  wire  pte_temp_flag_d = _GEN_5575[7]; // @[playground/src/cache/DCache.scala 649:102]
  wire [19:0] pte_temp_ppn = _GEN_5575[29:10]; // @[playground/src/cache/DCache.scala 649:102]
  wire  _T_57 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w; // @[playground/src/cache/DCache.scala 650:33]
  wire [1:0] _vpn_index_T_1 = vpn_index - 2'h1; // @[playground/src/cache/DCache.scala 659:38]
  wire [19:0] _GEN_5580 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_ppn : pte_ppn; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5582 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_d : pte_flag_d; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5583 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_a : pte_flag_a; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5584 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_g : pte_flag_g; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5585 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_u : pte_flag_u; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5586 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_x : pte_flag_x; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5587 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_w : pte_flag_w; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5588 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_r : pte_flag_r; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire  _GEN_5589 = pte_temp_flag_r | pte_temp_flag_x ? pte_temp_flag_v : pte_flag_v; // @[playground/src/cache/DCache.scala 653:54 655:25 569:28]
  wire [2:0] _GEN_5590 = pte_temp_flag_r | pte_temp_flag_x ? 3'h4 : 3'h1; // @[playground/src/cache/DCache.scala 653:54 656:25]
  wire [1:0] _GEN_5591 = pte_temp_flag_r | pte_temp_flag_x ? vpn_index : _vpn_index_T_1; // @[playground/src/cache/DCache.scala 568:28 653:54 659:25]
  wire [19:0] _GEN_5593 = pte_temp_flag_r | pte_temp_flag_x ? ppn : pte_temp_ppn; // @[playground/src/cache/DCache.scala 567:28 653:54]
  wire [2:0] _GEN_5595 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? 3'h0 : _GEN_5590; // @[playground/src/cache/DCache.scala 581:40 650:73]
  wire [19:0] _GEN_5597 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_ppn : _GEN_5580; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5599 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_d : _GEN_5582; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5600 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_a : _GEN_5583; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5601 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_g : _GEN_5584; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5602 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_u : _GEN_5585; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5603 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_x : _GEN_5586; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5604 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_w : _GEN_5587; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5605 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_r : _GEN_5588; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire  _GEN_5606 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? pte_flag_v : _GEN_5589; // @[playground/src/cache/DCache.scala 569:28 650:73]
  wire [1:0] _GEN_5607 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? vpn_index : _GEN_5591; // @[playground/src/cache/DCache.scala 568:28 650:73]
  wire [19:0] _GEN_5608 = ~pte_temp_flag_v | ~pte_temp_flag_r & pte_temp_flag_w ? ppn : _GEN_5593; // @[playground/src/cache/DCache.scala 567:28 650:73]
  wire  _GEN_5609 = cache_hit & _T_57; // @[playground/src/cache/DCache.scala 648:25 571:40]
  wire [2:0] _GEN_5610 = cache_hit ? _GEN_5595 : ptw_state; // @[playground/src/cache/DCache.scala 648:25 94:103]
  wire [19:0] _GEN_5612 = cache_hit ? _GEN_5597 : pte_ppn; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5614 = cache_hit ? _GEN_5599 : pte_flag_d; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5615 = cache_hit ? _GEN_5600 : pte_flag_a; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5616 = cache_hit ? _GEN_5601 : pte_flag_g; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5617 = cache_hit ? _GEN_5602 : pte_flag_u; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5618 = cache_hit ? _GEN_5603 : pte_flag_x; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5619 = cache_hit ? _GEN_5604 : pte_flag_w; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5620 = cache_hit ? _GEN_5605 : pte_flag_r; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire  _GEN_5621 = cache_hit ? _GEN_5606 : pte_flag_v; // @[playground/src/cache/DCache.scala 648:25 569:28]
  wire [1:0] _GEN_5622 = cache_hit ? _GEN_5607 : vpn_index; // @[playground/src/cache/DCache.scala 648:25 568:28]
  wire [19:0] _GEN_5623 = cache_hit ? _GEN_5608 : ppn; // @[playground/src/cache/DCache.scala 648:25 567:28]
  wire  _GEN_5624 = cache_hit ? _GEN_5405 : 1'h1; // @[playground/src/cache/DCache.scala 648:25 669:31]
  wire [2:0] _GEN_5625 = cache_hit ? _GEN_5056 : 3'h3; // @[playground/src/cache/DCache.scala 648:25 670:31]
  wire  _GEN_5626 = ~ptw_scratch_replace & _GEN_5609; // @[playground/src/cache/DCache.scala 647:34 571:40]
  wire [2:0] _GEN_5627 = ~ptw_scratch_replace ? _GEN_5610 : ptw_state; // @[playground/src/cache/DCache.scala 647:34 94:103]
  wire [19:0] _GEN_5629 = ~ptw_scratch_replace ? _GEN_5612 : pte_ppn; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5631 = ~ptw_scratch_replace ? _GEN_5614 : pte_flag_d; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5632 = ~ptw_scratch_replace ? _GEN_5615 : pte_flag_a; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5633 = ~ptw_scratch_replace ? _GEN_5616 : pte_flag_g; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5634 = ~ptw_scratch_replace ? _GEN_5617 : pte_flag_u; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5635 = ~ptw_scratch_replace ? _GEN_5618 : pte_flag_x; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5636 = ~ptw_scratch_replace ? _GEN_5619 : pte_flag_w; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5637 = ~ptw_scratch_replace ? _GEN_5620 : pte_flag_r; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire  _GEN_5638 = ~ptw_scratch_replace ? _GEN_5621 : pte_flag_v; // @[playground/src/cache/DCache.scala 569:28 647:34]
  wire [1:0] _GEN_5639 = ~ptw_scratch_replace ? _GEN_5622 : vpn_index; // @[playground/src/cache/DCache.scala 568:28 647:34]
  wire [19:0] _GEN_5640 = ~ptw_scratch_replace ? _GEN_5623 : ppn; // @[playground/src/cache/DCache.scala 567:28 647:34]
  wire  _GEN_5641 = ~ptw_scratch_replace ? _GEN_5624 : _GEN_5405; // @[playground/src/cache/DCache.scala 647:34]
  wire [2:0] _GEN_5642 = ~ptw_scratch_replace ? _GEN_5625 : _GEN_5056; // @[playground/src/cache/DCache.scala 647:34]
  wire  _GEN_5643 = _T_34 ? 1'h0 : _GEN_5065; // @[playground/src/cache/DCache.scala 675:28 676:17]
  wire  pte_temp_1_flag_v = io_axi_r_bits_data[0]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_r = io_axi_r_bits_data[1]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_w = io_axi_r_bits_data[2]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_x = io_axi_r_bits_data[3]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_u = io_axi_r_bits_data[4]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_g = io_axi_r_bits_data[5]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_a = io_axi_r_bits_data[6]; // @[playground/src/cache/DCache.scala 680:51]
  wire  pte_temp_1_flag_d = io_axi_r_bits_data[7]; // @[playground/src/cache/DCache.scala 680:51]
  wire [19:0] pte_temp_1_ppn = io_axi_r_bits_data[29:10]; // @[playground/src/cache/DCache.scala 680:51]
  wire  _T_68 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w; // @[playground/src/cache/DCache.scala 681:31]
  wire [19:0] _GEN_5648 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_ppn : pte_ppn; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5650 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_d : pte_flag_d; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5651 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_a : pte_flag_a; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5652 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_g : pte_flag_g; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5653 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_u : pte_flag_u; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5654 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_x : pte_flag_x; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5655 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_w : pte_flag_w; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5656 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_r : pte_flag_r; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire  _GEN_5657 = pte_temp_1_flag_r | pte_temp_1_flag_x ? pte_temp_1_flag_v : pte_flag_v; // @[playground/src/cache/DCache.scala 684:52 686:23 569:28]
  wire [2:0] _GEN_5658 = pte_temp_1_flag_r | pte_temp_1_flag_x ? 3'h4 : 3'h1; // @[playground/src/cache/DCache.scala 684:52 687:23]
  wire [1:0] _GEN_5659 = pte_temp_1_flag_r | pte_temp_1_flag_x ? vpn_index : _vpn_index_T_1; // @[playground/src/cache/DCache.scala 568:28 684:52 690:23]
  wire [19:0] _GEN_5661 = pte_temp_1_flag_r | pte_temp_1_flag_x ? ppn : pte_temp_1_ppn; // @[playground/src/cache/DCache.scala 567:28 684:52]
  wire [2:0] _GEN_5663 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? 3'h0 : _GEN_5658; // @[playground/src/cache/DCache.scala 581:40 681:71]
  wire [19:0] _GEN_5665 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_ppn : _GEN_5648; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5667 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_d : _GEN_5650; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5668 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_a : _GEN_5651; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5669 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_g : _GEN_5652; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5670 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_u : _GEN_5653; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5671 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_x : _GEN_5654; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5672 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_w : _GEN_5655; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5673 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_r : _GEN_5656; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire  _GEN_5674 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? pte_flag_v : _GEN_5657; // @[playground/src/cache/DCache.scala 569:28 681:71]
  wire [1:0] _GEN_5675 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? vpn_index : _GEN_5659; // @[playground/src/cache/DCache.scala 568:28 681:71]
  wire [19:0] _GEN_5676 = ~pte_temp_1_flag_v | ~pte_temp_1_flag_r & pte_temp_1_flag_w ? ppn : _GEN_5661; // @[playground/src/cache/DCache.scala 567:28 681:71]
  wire  _GEN_5677 = _T_18 ? 1'h0 : _GEN_5066; // @[playground/src/cache/DCache.scala 678:27 679:16]
  wire  _GEN_5678 = _T_18 & _T_68; // @[playground/src/cache/DCache.scala 678:27 571:40]
  wire [2:0] _GEN_5679 = _T_18 ? _GEN_5663 : ptw_state; // @[playground/src/cache/DCache.scala 678:27 94:103]
  wire [19:0] _GEN_5681 = _T_18 ? _GEN_5665 : pte_ppn; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5683 = _T_18 ? _GEN_5667 : pte_flag_d; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5684 = _T_18 ? _GEN_5668 : pte_flag_a; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5685 = _T_18 ? _GEN_5669 : pte_flag_g; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5686 = _T_18 ? _GEN_5670 : pte_flag_u; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5687 = _T_18 ? _GEN_5671 : pte_flag_x; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5688 = _T_18 ? _GEN_5672 : pte_flag_w; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5689 = _T_18 ? _GEN_5673 : pte_flag_r; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire  _GEN_5690 = _T_18 ? _GEN_5674 : pte_flag_v; // @[playground/src/cache/DCache.scala 678:27 569:28]
  wire [1:0] _GEN_5691 = _T_18 ? _GEN_5675 : vpn_index; // @[playground/src/cache/DCache.scala 678:27 568:28]
  wire [19:0] _GEN_5692 = _T_18 ? _GEN_5676 : ppn; // @[playground/src/cache/DCache.scala 678:27 567:28]
  wire  _T_75 = ~pte_flag_r; // @[playground/src/cache/DCache.scala 706:18]
  wire  _T_76 = ~pte_flag_x; // @[playground/src/cache/DCache.scala 706:33]
  wire  _T_80 = pte_flag_u & ~mstatus_sum; // @[playground/src/cache/DCache.scala 587:25]
  wire [2:0] _GEN_5694 = pte_flag_u & ~mstatus_sum ? 3'h0 : 3'h5; // @[playground/src/cache/DCache.scala 587:34 581:40 590:21]
  wire  _T_82 = ~pte_flag_u; // @[playground/src/cache/DCache.scala 594:14]
  wire [2:0] _GEN_5696 = ~pte_flag_u ? 3'h0 : 3'h5; // @[playground/src/cache/DCache.scala 594:27 581:40 597:21]
  wire  _GEN_5697 = 2'h0 == mode & _T_82; // @[playground/src/cache/DCache.scala 585:18 571:40]
  wire [2:0] _GEN_5698 = 2'h0 == mode ? _GEN_5696 : ptw_state; // @[playground/src/cache/DCache.scala 585:18 94:103]
  wire  _GEN_5699 = 2'h1 == mode ? _T_80 : _GEN_5697; // @[playground/src/cache/DCache.scala 585:18]
  wire [2:0] _GEN_5700 = 2'h1 == mode ? _GEN_5694 : _GEN_5698; // @[playground/src/cache/DCache.scala 585:18]
  wire  _GEN_5701 = ~pte_flag_r & ~pte_flag_x | _GEN_5699; // @[playground/src/cache/DCache.scala 579:40 706:46]
  wire [2:0] _GEN_5702 = ~pte_flag_r & ~pte_flag_x ? 3'h0 : _GEN_5700; // @[playground/src/cache/DCache.scala 581:40 706:46]
  wire  _GEN_5711 = _T_75 | _GEN_5699; // @[playground/src/cache/DCache.scala 712:31 579:40]
  wire [2:0] _GEN_5712 = _T_75 ? 3'h0 : _GEN_5700; // @[playground/src/cache/DCache.scala 712:31 581:40]
  wire  _GEN_5713 = mstatus_mxr ? _GEN_5701 : _GEN_5711; // @[playground/src/cache/DCache.scala 705:21]
  wire [2:0] _GEN_5714 = mstatus_mxr ? _GEN_5702 : _GEN_5712; // @[playground/src/cache/DCache.scala 705:21]
  wire  _GEN_5723 = ~pte_flag_w | _GEN_5699; // @[playground/src/cache/DCache.scala 720:29 579:40]
  wire [2:0] _GEN_5724 = ~pte_flag_w ? 3'h0 : _GEN_5700; // @[playground/src/cache/DCache.scala 720:29 581:40]
  wire  _GEN_5733 = _T_76 | _GEN_5699; // @[playground/src/cache/DCache.scala 727:29 579:40]
  wire [2:0] _GEN_5734 = _T_76 ? 3'h0 : _GEN_5700; // @[playground/src/cache/DCache.scala 727:29 581:40]
  wire  _GEN_5735 = 2'h0 == io_cpu_tlb_ptw_access_type & _GEN_5733; // @[playground/src/cache/DCache.scala 703:27 571:40]
  wire [2:0] _GEN_5736 = 2'h0 == io_cpu_tlb_ptw_access_type ? _GEN_5734 : ptw_state; // @[playground/src/cache/DCache.scala 703:27 94:103]
  wire  _GEN_5737 = 2'h2 == io_cpu_tlb_ptw_access_type ? _GEN_5723 : _GEN_5735; // @[playground/src/cache/DCache.scala 703:27]
  wire [2:0] _GEN_5738 = 2'h2 == io_cpu_tlb_ptw_access_type ? _GEN_5724 : _GEN_5736; // @[playground/src/cache/DCache.scala 703:27]
  wire  _GEN_5739 = 2'h1 == io_cpu_tlb_ptw_access_type ? _GEN_5713 : _GEN_5737; // @[playground/src/cache/DCache.scala 703:27]
  wire [2:0] _GEN_5740 = 2'h1 == io_cpu_tlb_ptw_access_type ? _GEN_5714 : _GEN_5738; // @[playground/src/cache/DCache.scala 703:27]
  wire  _T_109 = |pte_ppn[8:0]; // @[playground/src/cache/DCache.scala 738:65]
  wire  _T_121 = _vpnn_T_2 & (|pte_ppn[17:9] | _T_109); // @[playground/src/cache/DCache.scala 739:31]
  wire  _T_122 = _vpnn_T_1 & |pte_ppn[8:0] | _T_121; // @[playground/src/cache/DCache.scala 738:69]
  wire  _T_123 = vpn_index > 2'h0 & _T_122; // @[playground/src/cache/DCache.scala 737:25]
  wire  _T_128 = ~pte_flag_a | io_cpu_tlb_ptw_access_type == 2'h2 & ~pte_flag_d; // @[playground/src/cache/DCache.scala 743:30]
  wire [1:0] _GEN_5741 = _vpnn_T_1 ? pte_ppn[19:18] : pte_ppn[19:18]; // @[playground/src/cache/DCache.scala 757:39 758:24 763:19]
  wire [8:0] _GEN_5742 = _vpnn_T_1 ? pte_ppn[17:9] : pte_ppn[17:9]; // @[playground/src/cache/DCache.scala 757:39 759:24 763:19]
  wire [8:0] _GEN_5743 = _vpnn_T_1 ? vpn_vpn0 : pte_ppn[8:0]; // @[playground/src/cache/DCache.scala 757:39 760:24 763:19]
  wire [17:0] _GEN_5744 = _vpnn_T_1 ? 18'h3fe00 : 18'h3ffff; // @[playground/src/cache/DCache.scala 757:39 761:24 747:29]
  wire [1:0] ppn_set_ppn2 = _vpnn_T_2 ? pte_ppn[19:18] : _GEN_5741; // @[playground/src/cache/DCache.scala 752:33 753:24]
  wire [8:0] ppn_set_ppn1 = _vpnn_T_2 ? vpn_vpn1 : _GEN_5742; // @[playground/src/cache/DCache.scala 752:33 754:24]
  wire [8:0] ppn_set_ppn0 = _vpnn_T_2 ? vpn_vpn0 : _GEN_5743; // @[playground/src/cache/DCache.scala 752:33 755:24]
  wire [10:0] io_cpu_tlb_ptw_pte_bits_entry_ppn_hi = {ppn_set_ppn2,ppn_set_ppn1}; // @[playground/src/cache/DCache.scala 765:54]
  wire  _GEN_5765 = _T_123 | _T_128; // @[playground/src/cache/DCache.scala 580:40 741:9]
  wire  _GEN_5780 = 3'h5 == ptw_state & _GEN_5765; // @[playground/src/cache/DCache.scala 603:21 574:40]
  wire [2:0] _GEN_5781 = 3'h5 == ptw_state ? 3'h0 : ptw_state; // @[playground/src/cache/DCache.scala 603:21 94:103]
  wire  _GEN_5794 = 3'h4 == ptw_state ? _GEN_5739 : 3'h5 == ptw_state; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5795 = 3'h4 == ptw_state ? _GEN_5739 : _GEN_5780; // @[playground/src/cache/DCache.scala 603:21]
  wire [2:0] _GEN_5796 = 3'h4 == ptw_state ? _GEN_5740 : _GEN_5781; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5809 = 3'h3 == ptw_state ? _GEN_5643 : _GEN_5065; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5810 = 3'h3 == ptw_state ? _GEN_5677 : _GEN_5066; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5811 = 3'h3 == ptw_state ? _GEN_5678 : _GEN_5794; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5812 = 3'h3 == ptw_state ? _GEN_5678 : _GEN_5795; // @[playground/src/cache/DCache.scala 603:21]
  wire [2:0] _GEN_5813 = 3'h3 == ptw_state ? _GEN_5679 : _GEN_5796; // @[playground/src/cache/DCache.scala 603:21]
  wire [19:0] _GEN_5815 = 3'h3 == ptw_state ? _GEN_5681 : pte_ppn; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5817 = 3'h3 == ptw_state ? _GEN_5683 : pte_flag_d; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5818 = 3'h3 == ptw_state ? _GEN_5684 : pte_flag_a; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5819 = 3'h3 == ptw_state ? _GEN_5685 : pte_flag_g; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5820 = 3'h3 == ptw_state ? _GEN_5686 : pte_flag_u; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5821 = 3'h3 == ptw_state ? _GEN_5687 : pte_flag_x; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5822 = 3'h3 == ptw_state ? _GEN_5688 : pte_flag_w; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5823 = 3'h3 == ptw_state ? _GEN_5689 : pte_flag_r; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire  _GEN_5824 = 3'h3 == ptw_state ? _GEN_5690 : pte_flag_v; // @[playground/src/cache/DCache.scala 603:21 569:28]
  wire [1:0] _GEN_5825 = 3'h3 == ptw_state ? _GEN_5691 : vpn_index; // @[playground/src/cache/DCache.scala 603:21 568:28]
  wire [19:0] _GEN_5826 = 3'h3 == ptw_state ? _GEN_5692 : ppn; // @[playground/src/cache/DCache.scala 603:21 567:28]
  wire [5:0] _GEN_5839 = 3'h2 == ptw_state ? ptw_scratch_paddr_index : _bank_raddr_T_2; // @[playground/src/cache/DCache.scala 218:14 603:21 639:29]
  wire  _GEN_5844 = 3'h2 == ptw_state ? _GEN_5626 : _GEN_5811; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5845 = 3'h2 == ptw_state ? _GEN_5626 : _GEN_5812; // @[playground/src/cache/DCache.scala 603:21]
  wire [7:0] _GEN_5878 = 3'h1 == ptw_state ? _GEN_5421 : _GEN_5064; // @[playground/src/cache/DCache.scala 603:21]
  wire [5:0] _GEN_5882 = 3'h1 == ptw_state ? _GEN_5425 : _GEN_5839; // @[playground/src/cache/DCache.scala 603:21]
  wire  _GEN_5891 = 3'h1 == ptw_state ? 1'h0 : _GEN_5844; // @[playground/src/cache/DCache.scala 603:21 571:40]
  wire  _GEN_5892 = 3'h1 == ptw_state ? 1'h0 : _GEN_5845; // @[playground/src/cache/DCache.scala 603:21 574:40]
  wire [7:0] _GEN_5924 = 3'h0 == ptw_state ? _GEN_5064 : _GEN_5878; // @[playground/src/cache/DCache.scala 603:21]
  wire [7:0] _GEN_7927 = reset ? 8'h0 : _GEN_5924; // @[playground/src/cache/DCache.scala 259:{24,24}]
  wire [63:0] _GEN_7928 = reset ? 64'h0 : _GEN_5268; // @[playground/src/cache/DCache.scala 265:{24,24}]
  Queue writeFifo ( // @[playground/src/cache/DCache.scala 151:34]
    .clock(writeFifo_clock),
    .reset(writeFifo_reset),
    .io_enq_ready(writeFifo_io_enq_ready),
    .io_enq_valid(writeFifo_io_enq_valid),
    .io_enq_bits_data(writeFifo_io_enq_bits_data),
    .io_enq_bits_addr(writeFifo_io_enq_bits_addr),
    .io_enq_bits_strb(writeFifo_io_enq_bits_strb),
    .io_enq_bits_size(writeFifo_io_enq_bits_size),
    .io_deq_ready(writeFifo_io_deq_ready),
    .io_deq_valid(writeFifo_io_deq_valid),
    .io_deq_bits_data(writeFifo_io_deq_bits_data),
    .io_deq_bits_addr(writeFifo_io_deq_bits_addr),
    .io_deq_bits_strb(writeFifo_io_deq_bits_strb),
    .io_deq_bits_size(writeFifo_io_deq_bits_size)
  );
  LUTRam tagRam_0 ( // @[playground/src/cache/DCache.scala 226:37]
    .clock(tagRam_0_clock),
    .reset(tagRam_0_reset),
    .io_raddr(tagRam_0_io_raddr),
    .io_rdata(tagRam_0_io_rdata),
    .io_waddr(tagRam_0_io_waddr),
    .io_wdata(tagRam_0_io_wdata),
    .io_wen(tagRam_0_io_wen)
  );
  LUTRam tagRam_1 ( // @[playground/src/cache/DCache.scala 226:37]
    .clock(tagRam_1_clock),
    .reset(tagRam_1_reset),
    .io_raddr(tagRam_1_io_raddr),
    .io_rdata(tagRam_1_io_rdata),
    .io_waddr(tagRam_1_io_waddr),
    .io_wdata(tagRam_1_io_wdata),
    .io_wen(tagRam_1_io_wen)
  );
  SimpleDualPortRam_16 bank_0 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_0_clock),
    .reset(bank_0_reset),
    .io_raddr(bank_0_io_raddr),
    .io_rdata(bank_0_io_rdata),
    .io_waddr(bank_0_io_waddr),
    .io_wen(bank_0_io_wen),
    .io_wstrb(bank_0_io_wstrb),
    .io_wdata(bank_0_io_wdata)
  );
  SimpleDualPortRam_16 bank_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_1_clock),
    .reset(bank_1_reset),
    .io_raddr(bank_1_io_raddr),
    .io_rdata(bank_1_io_rdata),
    .io_waddr(bank_1_io_waddr),
    .io_wen(bank_1_io_wen),
    .io_wstrb(bank_1_io_wstrb),
    .io_wdata(bank_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_2 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_2_clock),
    .reset(bank_2_reset),
    .io_raddr(bank_2_io_raddr),
    .io_rdata(bank_2_io_rdata),
    .io_waddr(bank_2_io_waddr),
    .io_wen(bank_2_io_wen),
    .io_wstrb(bank_2_io_wstrb),
    .io_wdata(bank_2_io_wdata)
  );
  SimpleDualPortRam_16 bank_3 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_3_clock),
    .reset(bank_3_reset),
    .io_raddr(bank_3_io_raddr),
    .io_rdata(bank_3_io_rdata),
    .io_waddr(bank_3_io_waddr),
    .io_wen(bank_3_io_wen),
    .io_wstrb(bank_3_io_wstrb),
    .io_wdata(bank_3_io_wdata)
  );
  SimpleDualPortRam_16 bank_4 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_4_clock),
    .reset(bank_4_reset),
    .io_raddr(bank_4_io_raddr),
    .io_rdata(bank_4_io_rdata),
    .io_waddr(bank_4_io_waddr),
    .io_wen(bank_4_io_wen),
    .io_wstrb(bank_4_io_wstrb),
    .io_wdata(bank_4_io_wdata)
  );
  SimpleDualPortRam_16 bank_5 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_5_clock),
    .reset(bank_5_reset),
    .io_raddr(bank_5_io_raddr),
    .io_rdata(bank_5_io_rdata),
    .io_waddr(bank_5_io_waddr),
    .io_wen(bank_5_io_wen),
    .io_wstrb(bank_5_io_wstrb),
    .io_wdata(bank_5_io_wdata)
  );
  SimpleDualPortRam_16 bank_6 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_6_clock),
    .reset(bank_6_reset),
    .io_raddr(bank_6_io_raddr),
    .io_rdata(bank_6_io_rdata),
    .io_waddr(bank_6_io_waddr),
    .io_wen(bank_6_io_wen),
    .io_wstrb(bank_6_io_wstrb),
    .io_wdata(bank_6_io_wdata)
  );
  SimpleDualPortRam_16 bank_7 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_7_clock),
    .reset(bank_7_reset),
    .io_raddr(bank_7_io_raddr),
    .io_rdata(bank_7_io_rdata),
    .io_waddr(bank_7_io_waddr),
    .io_wen(bank_7_io_wen),
    .io_wstrb(bank_7_io_wstrb),
    .io_wdata(bank_7_io_wdata)
  );
  SimpleDualPortRam_16 bank_0_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_0_1_clock),
    .reset(bank_0_1_reset),
    .io_raddr(bank_0_1_io_raddr),
    .io_rdata(bank_0_1_io_rdata),
    .io_waddr(bank_0_1_io_waddr),
    .io_wen(bank_0_1_io_wen),
    .io_wstrb(bank_0_1_io_wstrb),
    .io_wdata(bank_0_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_1_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_1_1_clock),
    .reset(bank_1_1_reset),
    .io_raddr(bank_1_1_io_raddr),
    .io_rdata(bank_1_1_io_rdata),
    .io_waddr(bank_1_1_io_waddr),
    .io_wen(bank_1_1_io_wen),
    .io_wstrb(bank_1_1_io_wstrb),
    .io_wdata(bank_1_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_2_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_2_1_clock),
    .reset(bank_2_1_reset),
    .io_raddr(bank_2_1_io_raddr),
    .io_rdata(bank_2_1_io_rdata),
    .io_waddr(bank_2_1_io_waddr),
    .io_wen(bank_2_1_io_wen),
    .io_wstrb(bank_2_1_io_wstrb),
    .io_wdata(bank_2_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_3_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_3_1_clock),
    .reset(bank_3_1_reset),
    .io_raddr(bank_3_1_io_raddr),
    .io_rdata(bank_3_1_io_rdata),
    .io_waddr(bank_3_1_io_waddr),
    .io_wen(bank_3_1_io_wen),
    .io_wstrb(bank_3_1_io_wstrb),
    .io_wdata(bank_3_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_4_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_4_1_clock),
    .reset(bank_4_1_reset),
    .io_raddr(bank_4_1_io_raddr),
    .io_rdata(bank_4_1_io_rdata),
    .io_waddr(bank_4_1_io_waddr),
    .io_wen(bank_4_1_io_wen),
    .io_wstrb(bank_4_1_io_wstrb),
    .io_wdata(bank_4_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_5_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_5_1_clock),
    .reset(bank_5_1_reset),
    .io_raddr(bank_5_1_io_raddr),
    .io_rdata(bank_5_1_io_rdata),
    .io_waddr(bank_5_1_io_waddr),
    .io_wen(bank_5_1_io_wen),
    .io_wstrb(bank_5_1_io_wstrb),
    .io_wdata(bank_5_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_6_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_6_1_clock),
    .reset(bank_6_1_reset),
    .io_raddr(bank_6_1_io_raddr),
    .io_rdata(bank_6_1_io_rdata),
    .io_waddr(bank_6_1_io_waddr),
    .io_wen(bank_6_1_io_wen),
    .io_wstrb(bank_6_1_io_wstrb),
    .io_wdata(bank_6_1_io_wdata)
  );
  SimpleDualPortRam_16 bank_7_1 ( // @[playground/src/cache/DCache.scala 228:38]
    .clock(bank_7_1_clock),
    .reset(bank_7_1_reset),
    .io_raddr(bank_7_1_io_raddr),
    .io_rdata(bank_7_1_io_rdata),
    .io_waddr(bank_7_1_io_waddr),
    .io_wen(bank_7_1_io_wen),
    .io_wstrb(bank_7_1_io_wstrb),
    .io_wdata(bank_7_1_io_wdata)
  );
  assign io_cpu_rdata = _use_next_addr_T_1 ? saved_rdata : _GEN_15; // @[playground/src/cache/DCache.scala 211:22]
  assign io_cpu_access_fault = access_fault; // @[playground/src/cache/DCache.scala 286:23]
  assign io_cpu_page_fault = page_fault; // @[playground/src/cache/DCache.scala 287:23]
  assign io_cpu_dcache_ready = ~dcache_stall; // @[playground/src/cache/DCache.scala 207:26]
  assign io_cpu_tlb_en = io_cpu_en; // @[playground/src/cache/DCache.scala 215:26]
  assign io_cpu_tlb_vaddr = io_cpu_addr; // @[playground/src/cache/DCache.scala 213:26]
  assign io_cpu_tlb_complete_single_request = io_cpu_complete_single_request; // @[playground/src/cache/DCache.scala 575:40]
  assign io_cpu_tlb_access_type = io_cpu_en & _mmio_read_stall_T ? 2'h2 : 2'h1; // @[playground/src/cache/DCache.scala 214:32]
  assign io_cpu_tlb_ptw_vpn_ready = 3'h0 == state ? _GEN_1858 : _GEN_5052; // @[playground/src/cache/DCache.scala 316:17]
  assign io_cpu_tlb_ptw_pte_valid = 3'h0 == ptw_state ? 1'h0 : _GEN_5891; // @[playground/src/cache/DCache.scala 603:21 571:40]
  assign io_cpu_tlb_ptw_pte_bits_access_fault = 1'h0; // @[playground/src/cache/DCache.scala 573:40]
  assign io_cpu_tlb_ptw_pte_bits_page_fault = 3'h0 == ptw_state ? 1'h0 : _GEN_5892; // @[playground/src/cache/DCache.scala 603:21 574:40]
  assign io_cpu_tlb_ptw_pte_bits_entry_ppn = {io_cpu_tlb_ptw_pte_bits_entry_ppn_hi,ppn_set_ppn0}; // @[playground/src/cache/DCache.scala 765:54]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_d = pte_flag_d; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_g = pte_flag_g; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_u = pte_flag_u; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_x = pte_flag_x; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_w = pte_flag_w; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_r = pte_flag_r; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_entry_flag_v = pte_flag_v; // @[playground/src/cache/DCache.scala 743:82 750:39]
  assign io_cpu_tlb_ptw_pte_bits_rmask = _vpnn_T_2 ? 18'h0 : _GEN_5744; // @[playground/src/cache/DCache.scala 752:33 756:24]
  assign io_axi_ar_valid = arvalid; // @[playground/src/cache/DCache.scala 262:19]
  assign io_axi_ar_bits_addr = ar_addr; // @[playground/src/cache/DCache.scala 261:18]
  assign io_axi_ar_bits_len = ar_len; // @[playground/src/cache/DCache.scala 261:18]
  assign io_axi_ar_bits_size = ar_size; // @[playground/src/cache/DCache.scala 261:18]
  assign io_axi_r_ready = rready; // @[playground/src/cache/DCache.scala 264:18]
  assign io_axi_aw_valid = awvalid; // @[playground/src/cache/DCache.scala 268:19]
  assign io_axi_aw_bits_addr = aw_addr; // @[playground/src/cache/DCache.scala 267:18]
  assign io_axi_aw_bits_len = aw_len; // @[playground/src/cache/DCache.scala 267:18]
  assign io_axi_aw_bits_size = aw_size; // @[playground/src/cache/DCache.scala 267:18]
  assign io_axi_w_valid = wvalid; // @[playground/src/cache/DCache.scala 273:22]
  assign io_axi_w_bits_data = w_data; // @[playground/src/cache/DCache.scala 271:17]
  assign io_axi_w_bits_strb = w_strb; // @[playground/src/cache/DCache.scala 271:17]
  assign io_axi_w_bits_last = w_last & wvalid; // @[playground/src/cache/DCache.scala 272:32]
  assign io_axi_b_ready = 1'h1; // @[playground/src/cache/DCache.scala 275:18]
  assign writeFifo_clock = clock;
  assign writeFifo_reset = reset;
  assign writeFifo_io_enq_valid = 3'h0 == state & _GEN_1655; // @[playground/src/cache/DCache.scala 316:17 155:26]
  assign writeFifo_io_enq_bits_data = 3'h0 == state ? _GEN_1659 : 64'h0; // @[playground/src/cache/DCache.scala 316:17 156:26]
  assign writeFifo_io_enq_bits_addr = 3'h0 == state ? _GEN_1656 : 64'h0; // @[playground/src/cache/DCache.scala 316:17 156:26]
  assign writeFifo_io_enq_bits_strb = 3'h0 == state ? _GEN_1658 : 8'h0; // @[playground/src/cache/DCache.scala 316:17 156:26]
  assign writeFifo_io_enq_bits_size = _GEN_5059[2:0];
  assign writeFifo_io_deq_ready = writeFifo_axi_busy ? 1'h0 : _GEN_280; // @[playground/src/cache/DCache.scala 157:26 290:28]
  assign tagRam_0_clock = clock;
  assign tagRam_0_reset = reset;
  assign tagRam_0_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 603:21 239:26]
  assign tagRam_0_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign tagRam_0_io_wdata = tag_wdata; // @[playground/src/cache/DCache.scala 244:26]
  assign tagRam_0_io_wen = tag_wstrb_0; // @[playground/src/cache/DCache.scala 242:26]
  assign tagRam_1_clock = clock;
  assign tagRam_1_reset = reset;
  assign tagRam_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 603:21 239:26]
  assign tagRam_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign tagRam_1_io_wdata = tag_wdata; // @[playground/src/cache/DCache.scala 244:26]
  assign tagRam_1_io_wen = tag_wstrb_1; // @[playground/src/cache/DCache.scala 242:26]
  assign bank_0_clock = clock;
  assign bank_0_reset = reset;
  assign bank_0_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_0_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_0_io_wen = |replace_wstrb_0_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_0_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_0_0 : _replace_wstrb_0_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_0_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_1_clock = clock;
  assign bank_1_reset = reset;
  assign bank_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_1_io_wen = |replace_wstrb_1_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_1_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_1_0 : _replace_wstrb_1_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_2_clock = clock;
  assign bank_2_reset = reset;
  assign bank_2_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_2_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_2_io_wen = |replace_wstrb_2_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_2_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_2_0 : _replace_wstrb_2_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_2_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_3_clock = clock;
  assign bank_3_reset = reset;
  assign bank_3_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_3_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_3_io_wen = |replace_wstrb_3_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_3_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_3_0 : _replace_wstrb_3_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_3_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_4_clock = clock;
  assign bank_4_reset = reset;
  assign bank_4_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_4_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_4_io_wen = |replace_wstrb_4_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_4_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_4_0 : _replace_wstrb_4_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_4_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_5_clock = clock;
  assign bank_5_reset = reset;
  assign bank_5_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_5_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_5_io_wen = |replace_wstrb_5_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_5_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_5_0 : _replace_wstrb_5_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_5_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_6_clock = clock;
  assign bank_6_reset = reset;
  assign bank_6_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_6_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_6_io_wen = |replace_wstrb_6_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_6_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_6_0 : _replace_wstrb_6_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_6_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_7_clock = clock;
  assign bank_7_reset = reset;
  assign bank_7_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_7_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_7_io_wen = |replace_wstrb_7_0; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_7_io_wstrb = _replace_wstrb_0_0_T_6 ? wstrb_7_0 : _replace_wstrb_7_0_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_7_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_0_1_clock = clock;
  assign bank_0_1_reset = reset;
  assign bank_0_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_0_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_0_1_io_wen = |replace_wstrb_0_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_0_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_0_1 : _replace_wstrb_0_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_0_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_1_1_clock = clock;
  assign bank_1_1_reset = reset;
  assign bank_1_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_1_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_1_1_io_wen = |replace_wstrb_1_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_1_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_1_1 : _replace_wstrb_1_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_1_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_2_1_clock = clock;
  assign bank_2_1_reset = reset;
  assign bank_2_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_2_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_2_1_io_wen = |replace_wstrb_2_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_2_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_2_1 : _replace_wstrb_2_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_2_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_3_1_clock = clock;
  assign bank_3_1_reset = reset;
  assign bank_3_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_3_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_3_1_io_wen = |replace_wstrb_3_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_3_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_3_1 : _replace_wstrb_3_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_3_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_4_1_clock = clock;
  assign bank_4_1_reset = reset;
  assign bank_4_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_4_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_4_1_io_wen = |replace_wstrb_4_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_4_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_4_1 : _replace_wstrb_4_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_4_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_5_1_clock = clock;
  assign bank_5_1_reset = reset;
  assign bank_5_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_5_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_5_1_io_wen = |replace_wstrb_5_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_5_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_5_1 : _replace_wstrb_5_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_5_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_6_1_clock = clock;
  assign bank_6_1_reset = reset;
  assign bank_6_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_6_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_6_1_io_wen = |replace_wstrb_6_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_6_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_6_1 : _replace_wstrb_6_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_6_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  assign bank_7_1_clock = clock;
  assign bank_7_1_reset = reset;
  assign bank_7_1_io_raddr = 3'h0 == ptw_state ? _bank_raddr_T_2 : _GEN_5882; // @[playground/src/cache/DCache.scala 218:14 603:21]
  assign bank_7_1_io_waddr = 3'h0 == ptw_state ? io_cpu_addr[11:6] : _GEN_5884; // @[playground/src/cache/DCache.scala 173:17 603:21]
  assign bank_7_1_io_wen = |replace_wstrb_7_1; // @[playground/src/cache/DCache.scala 234:47]
  assign bank_7_1_io_wstrb = _replace_wstrb_0_1_T_6 ? wstrb_7_1 : _replace_wstrb_7_1_T_9; // @[playground/src/cache/DCache.scala 251:33]
  assign bank_7_1_io_wdata = state == 3'h3 ? io_axi_r_bits_data : io_cpu_wdata; // @[playground/src/cache/DCache.scala 175:26]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/cache/DCache.scala 90:94]
      state <= 3'h0; // @[playground/src/cache/DCache.scala 90:94]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      state <= _GEN_5056;
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      state <= _GEN_5056;
    end else if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      state <= _GEN_5642;
    end else begin
      state <= _GEN_5056;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 94:103]
      ptw_state <= 3'h0; // @[playground/src/cache/DCache.scala 94:103]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      if (_T_50) begin // @[playground/src/cache/DCache.scala 606:37]
        ptw_state <= 3'h1; // @[playground/src/cache/DCache.scala 609:19]
      end
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      if (pte_uncached) begin // @[playground/src/cache/DCache.scala 622:26]
        ptw_state <= 3'h3; // @[playground/src/cache/DCache.scala 628:19]
      end else begin
        ptw_state <= 3'h2; // @[playground/src/cache/DCache.scala 633:31]
      end
    end else if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      ptw_state <= _GEN_5627;
    end else begin
      ptw_state <= _GEN_5813;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 101:28]
      ptw_scratch_paddr_tag <= 20'h0; // @[playground/src/cache/DCache.scala 101:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
        if (!(pte_uncached)) begin // @[playground/src/cache/DCache.scala 622:26]
          ptw_scratch_paddr_tag <= ptw_addr_tag; // @[playground/src/cache/DCache.scala 634:31]
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 101:28]
      ptw_scratch_paddr_index <= 6'h0; // @[playground/src/cache/DCache.scala 101:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
        if (!(pte_uncached)) begin // @[playground/src/cache/DCache.scala 622:26]
          ptw_scratch_paddr_index <= ptw_addr_index; // @[playground/src/cache/DCache.scala 634:31]
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 101:28]
      ptw_scratch_paddr_offset <= 6'h0; // @[playground/src/cache/DCache.scala 101:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
        if (!(pte_uncached)) begin // @[playground/src/cache/DCache.scala 622:26]
          ptw_scratch_paddr_offset <= ptw_addr_offset; // @[playground/src/cache/DCache.scala 634:31]
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 101:28]
      ptw_scratch_replace <= 1'h0; // @[playground/src/cache/DCache.scala 101:28]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      ptw_scratch_replace <= _GEN_5405;
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      ptw_scratch_replace <= _GEN_5431;
    end else if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      ptw_scratch_replace <= _GEN_5641;
    end else begin
      ptw_scratch_replace <= _GEN_5405;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 101:28]
      ptw_scratch_dcache_wait <= 1'h0; // @[playground/src/cache/DCache.scala 101:28]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          ptw_scratch_dcache_wait <= _GEN_4448;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_0_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_0_0 <= _GEN_4317;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_0_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_0_1 <= _GEN_4318;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_1_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_1_0 <= _GEN_4319;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_1_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_1_1 <= _GEN_4320;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_2_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_2_0 <= _GEN_4321;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_2_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_2_1 <= _GEN_4322;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_3_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_3_0 <= _GEN_4323;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_3_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_3_1 <= _GEN_4324;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_4_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_4_0 <= _GEN_4325;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_4_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_4_1 <= _GEN_4326;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_5_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_5_0 <= _GEN_4327;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_5_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_5_1 <= _GEN_4328;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_6_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_6_0 <= _GEN_4329;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_6_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_6_1 <= _GEN_4330;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_7_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_7_0 <= _GEN_4331;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_7_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_7_1 <= _GEN_4332;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_8_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_8_0 <= _GEN_4333;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_8_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_8_1 <= _GEN_4334;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_9_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_9_0 <= _GEN_4335;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_9_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_9_1 <= _GEN_4336;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_10_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_10_0 <= _GEN_4337;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_10_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_10_1 <= _GEN_4338;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_11_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_11_0 <= _GEN_4339;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_11_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_11_1 <= _GEN_4340;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_12_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_12_0 <= _GEN_4341;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_12_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_12_1 <= _GEN_4342;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_13_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_13_0 <= _GEN_4343;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_13_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_13_1 <= _GEN_4344;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_14_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_14_0 <= _GEN_4345;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_14_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_14_1 <= _GEN_4346;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_15_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_15_0 <= _GEN_4347;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_15_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_15_1 <= _GEN_4348;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_16_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_16_0 <= _GEN_4349;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_16_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_16_1 <= _GEN_4350;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_17_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_17_0 <= _GEN_4351;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_17_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_17_1 <= _GEN_4352;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_18_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_18_0 <= _GEN_4353;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_18_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_18_1 <= _GEN_4354;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_19_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_19_0 <= _GEN_4355;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_19_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_19_1 <= _GEN_4356;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_20_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_20_0 <= _GEN_4357;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_20_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_20_1 <= _GEN_4358;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_21_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_21_0 <= _GEN_4359;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_21_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_21_1 <= _GEN_4360;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_22_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_22_0 <= _GEN_4361;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_22_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_22_1 <= _GEN_4362;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_23_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_23_0 <= _GEN_4363;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_23_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_23_1 <= _GEN_4364;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_24_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_24_0 <= _GEN_4365;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_24_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_24_1 <= _GEN_4366;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_25_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_25_0 <= _GEN_4367;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_25_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_25_1 <= _GEN_4368;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_26_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_26_0 <= _GEN_4369;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_26_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_26_1 <= _GEN_4370;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_27_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_27_0 <= _GEN_4371;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_27_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_27_1 <= _GEN_4372;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_28_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_28_0 <= _GEN_4373;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_28_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_28_1 <= _GEN_4374;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_29_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_29_0 <= _GEN_4375;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_29_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_29_1 <= _GEN_4376;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_30_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_30_0 <= _GEN_4377;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_30_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_30_1 <= _GEN_4378;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_31_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_31_0 <= _GEN_4379;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_31_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_31_1 <= _GEN_4380;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_32_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_32_0 <= _GEN_4381;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_32_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_32_1 <= _GEN_4382;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_33_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_33_0 <= _GEN_4383;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_33_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_33_1 <= _GEN_4384;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_34_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_34_0 <= _GEN_4385;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_34_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_34_1 <= _GEN_4386;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_35_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_35_0 <= _GEN_4387;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_35_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_35_1 <= _GEN_4388;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_36_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_36_0 <= _GEN_4389;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_36_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_36_1 <= _GEN_4390;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_37_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_37_0 <= _GEN_4391;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_37_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_37_1 <= _GEN_4392;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_38_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_38_0 <= _GEN_4393;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_38_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_38_1 <= _GEN_4394;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_39_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_39_0 <= _GEN_4395;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_39_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_39_1 <= _GEN_4396;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_40_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_40_0 <= _GEN_4397;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_40_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_40_1 <= _GEN_4398;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_41_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_41_0 <= _GEN_4399;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_41_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_41_1 <= _GEN_4400;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_42_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_42_0 <= _GEN_4401;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_42_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_42_1 <= _GEN_4402;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_43_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_43_0 <= _GEN_4403;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_43_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_43_1 <= _GEN_4404;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_44_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_44_0 <= _GEN_4405;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_44_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_44_1 <= _GEN_4406;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_45_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_45_0 <= _GEN_4407;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_45_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_45_1 <= _GEN_4408;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_46_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_46_0 <= _GEN_4409;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_46_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_46_1 <= _GEN_4410;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_47_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_47_0 <= _GEN_4411;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_47_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_47_1 <= _GEN_4412;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_48_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_48_0 <= _GEN_4413;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_48_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_48_1 <= _GEN_4414;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_49_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_49_0 <= _GEN_4415;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_49_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_49_1 <= _GEN_4416;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_50_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_50_0 <= _GEN_4417;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_50_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_50_1 <= _GEN_4418;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_51_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_51_0 <= _GEN_4419;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_51_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_51_1 <= _GEN_4420;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_52_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_52_0 <= _GEN_4421;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_52_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_52_1 <= _GEN_4422;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_53_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_53_0 <= _GEN_4423;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_53_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_53_1 <= _GEN_4424;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_54_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_54_0 <= _GEN_4425;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_54_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_54_1 <= _GEN_4426;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_55_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_55_0 <= _GEN_4427;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_55_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_55_1 <= _GEN_4428;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_56_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_56_0 <= _GEN_4429;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_56_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_56_1 <= _GEN_4430;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_57_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_57_0 <= _GEN_4431;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_57_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_57_1 <= _GEN_4432;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_58_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_58_0 <= _GEN_4433;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_58_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_58_1 <= _GEN_4434;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_59_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_59_0 <= _GEN_4435;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_59_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_59_1 <= _GEN_4436;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_60_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_60_0 <= _GEN_4437;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_60_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_60_1 <= _GEN_4438;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_61_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_61_0 <= _GEN_4439;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_61_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_61_1 <= _GEN_4440;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_62_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_62_0 <= _GEN_4441;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_62_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_62_1 <= _GEN_4442;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_63_0 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_63_0 <= _GEN_4443;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 134:22]
      valid_63_1 <= 1'h0; // @[playground/src/cache/DCache.scala 134:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          valid_63_1 <= _GEN_4444;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_0_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_0_0 <= _GEN_1313;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_0_0 <= _GEN_2242;
      end else begin
        dirty_0_0 <= _GEN_4183;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_0_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_0_1 <= _GEN_1314;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_0_1 <= _GEN_2243;
      end else begin
        dirty_0_1 <= _GEN_4184;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_1_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_1_0 <= _GEN_1315;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_1_0 <= _GEN_2244;
      end else begin
        dirty_1_0 <= _GEN_4185;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_1_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_1_1 <= _GEN_1316;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_1_1 <= _GEN_2245;
      end else begin
        dirty_1_1 <= _GEN_4186;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_2_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_2_0 <= _GEN_1317;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_2_0 <= _GEN_2246;
      end else begin
        dirty_2_0 <= _GEN_4187;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_2_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_2_1 <= _GEN_1318;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_2_1 <= _GEN_2247;
      end else begin
        dirty_2_1 <= _GEN_4188;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_3_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_3_0 <= _GEN_1319;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_3_0 <= _GEN_2248;
      end else begin
        dirty_3_0 <= _GEN_4189;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_3_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_3_1 <= _GEN_1320;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_3_1 <= _GEN_2249;
      end else begin
        dirty_3_1 <= _GEN_4190;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_4_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_4_0 <= _GEN_1321;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_4_0 <= _GEN_2250;
      end else begin
        dirty_4_0 <= _GEN_4191;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_4_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_4_1 <= _GEN_1322;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_4_1 <= _GEN_2251;
      end else begin
        dirty_4_1 <= _GEN_4192;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_5_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_5_0 <= _GEN_1323;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_5_0 <= _GEN_2252;
      end else begin
        dirty_5_0 <= _GEN_4193;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_5_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_5_1 <= _GEN_1324;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_5_1 <= _GEN_2253;
      end else begin
        dirty_5_1 <= _GEN_4194;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_6_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_6_0 <= _GEN_1325;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_6_0 <= _GEN_2254;
      end else begin
        dirty_6_0 <= _GEN_4195;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_6_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_6_1 <= _GEN_1326;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_6_1 <= _GEN_2255;
      end else begin
        dirty_6_1 <= _GEN_4196;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_7_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_7_0 <= _GEN_1327;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_7_0 <= _GEN_2256;
      end else begin
        dirty_7_0 <= _GEN_4197;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_7_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_7_1 <= _GEN_1328;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_7_1 <= _GEN_2257;
      end else begin
        dirty_7_1 <= _GEN_4198;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_8_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_8_0 <= _GEN_1329;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_8_0 <= _GEN_2258;
      end else begin
        dirty_8_0 <= _GEN_4199;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_8_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_8_1 <= _GEN_1330;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_8_1 <= _GEN_2259;
      end else begin
        dirty_8_1 <= _GEN_4200;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_9_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_9_0 <= _GEN_1331;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_9_0 <= _GEN_2260;
      end else begin
        dirty_9_0 <= _GEN_4201;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_9_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_9_1 <= _GEN_1332;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_9_1 <= _GEN_2261;
      end else begin
        dirty_9_1 <= _GEN_4202;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_10_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_10_0 <= _GEN_1333;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_10_0 <= _GEN_2262;
      end else begin
        dirty_10_0 <= _GEN_4203;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_10_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_10_1 <= _GEN_1334;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_10_1 <= _GEN_2263;
      end else begin
        dirty_10_1 <= _GEN_4204;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_11_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_11_0 <= _GEN_1335;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_11_0 <= _GEN_2264;
      end else begin
        dirty_11_0 <= _GEN_4205;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_11_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_11_1 <= _GEN_1336;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_11_1 <= _GEN_2265;
      end else begin
        dirty_11_1 <= _GEN_4206;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_12_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_12_0 <= _GEN_1337;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_12_0 <= _GEN_2266;
      end else begin
        dirty_12_0 <= _GEN_4207;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_12_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_12_1 <= _GEN_1338;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_12_1 <= _GEN_2267;
      end else begin
        dirty_12_1 <= _GEN_4208;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_13_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_13_0 <= _GEN_1339;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_13_0 <= _GEN_2268;
      end else begin
        dirty_13_0 <= _GEN_4209;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_13_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_13_1 <= _GEN_1340;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_13_1 <= _GEN_2269;
      end else begin
        dirty_13_1 <= _GEN_4210;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_14_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_14_0 <= _GEN_1341;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_14_0 <= _GEN_2270;
      end else begin
        dirty_14_0 <= _GEN_4211;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_14_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_14_1 <= _GEN_1342;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_14_1 <= _GEN_2271;
      end else begin
        dirty_14_1 <= _GEN_4212;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_15_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_15_0 <= _GEN_1343;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_15_0 <= _GEN_2272;
      end else begin
        dirty_15_0 <= _GEN_4213;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_15_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_15_1 <= _GEN_1344;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_15_1 <= _GEN_2273;
      end else begin
        dirty_15_1 <= _GEN_4214;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_16_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_16_0 <= _GEN_1345;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_16_0 <= _GEN_2274;
      end else begin
        dirty_16_0 <= _GEN_4215;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_16_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_16_1 <= _GEN_1346;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_16_1 <= _GEN_2275;
      end else begin
        dirty_16_1 <= _GEN_4216;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_17_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_17_0 <= _GEN_1347;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_17_0 <= _GEN_2276;
      end else begin
        dirty_17_0 <= _GEN_4217;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_17_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_17_1 <= _GEN_1348;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_17_1 <= _GEN_2277;
      end else begin
        dirty_17_1 <= _GEN_4218;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_18_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_18_0 <= _GEN_1349;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_18_0 <= _GEN_2278;
      end else begin
        dirty_18_0 <= _GEN_4219;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_18_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_18_1 <= _GEN_1350;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_18_1 <= _GEN_2279;
      end else begin
        dirty_18_1 <= _GEN_4220;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_19_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_19_0 <= _GEN_1351;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_19_0 <= _GEN_2280;
      end else begin
        dirty_19_0 <= _GEN_4221;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_19_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_19_1 <= _GEN_1352;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_19_1 <= _GEN_2281;
      end else begin
        dirty_19_1 <= _GEN_4222;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_20_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_20_0 <= _GEN_1353;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_20_0 <= _GEN_2282;
      end else begin
        dirty_20_0 <= _GEN_4223;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_20_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_20_1 <= _GEN_1354;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_20_1 <= _GEN_2283;
      end else begin
        dirty_20_1 <= _GEN_4224;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_21_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_21_0 <= _GEN_1355;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_21_0 <= _GEN_2284;
      end else begin
        dirty_21_0 <= _GEN_4225;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_21_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_21_1 <= _GEN_1356;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_21_1 <= _GEN_2285;
      end else begin
        dirty_21_1 <= _GEN_4226;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_22_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_22_0 <= _GEN_1357;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_22_0 <= _GEN_2286;
      end else begin
        dirty_22_0 <= _GEN_4227;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_22_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_22_1 <= _GEN_1358;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_22_1 <= _GEN_2287;
      end else begin
        dirty_22_1 <= _GEN_4228;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_23_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_23_0 <= _GEN_1359;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_23_0 <= _GEN_2288;
      end else begin
        dirty_23_0 <= _GEN_4229;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_23_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_23_1 <= _GEN_1360;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_23_1 <= _GEN_2289;
      end else begin
        dirty_23_1 <= _GEN_4230;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_24_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_24_0 <= _GEN_1361;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_24_0 <= _GEN_2290;
      end else begin
        dirty_24_0 <= _GEN_4231;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_24_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_24_1 <= _GEN_1362;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_24_1 <= _GEN_2291;
      end else begin
        dirty_24_1 <= _GEN_4232;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_25_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_25_0 <= _GEN_1363;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_25_0 <= _GEN_2292;
      end else begin
        dirty_25_0 <= _GEN_4233;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_25_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_25_1 <= _GEN_1364;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_25_1 <= _GEN_2293;
      end else begin
        dirty_25_1 <= _GEN_4234;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_26_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_26_0 <= _GEN_1365;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_26_0 <= _GEN_2294;
      end else begin
        dirty_26_0 <= _GEN_4235;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_26_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_26_1 <= _GEN_1366;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_26_1 <= _GEN_2295;
      end else begin
        dirty_26_1 <= _GEN_4236;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_27_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_27_0 <= _GEN_1367;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_27_0 <= _GEN_2296;
      end else begin
        dirty_27_0 <= _GEN_4237;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_27_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_27_1 <= _GEN_1368;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_27_1 <= _GEN_2297;
      end else begin
        dirty_27_1 <= _GEN_4238;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_28_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_28_0 <= _GEN_1369;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_28_0 <= _GEN_2298;
      end else begin
        dirty_28_0 <= _GEN_4239;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_28_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_28_1 <= _GEN_1370;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_28_1 <= _GEN_2299;
      end else begin
        dirty_28_1 <= _GEN_4240;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_29_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_29_0 <= _GEN_1371;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_29_0 <= _GEN_2300;
      end else begin
        dirty_29_0 <= _GEN_4241;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_29_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_29_1 <= _GEN_1372;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_29_1 <= _GEN_2301;
      end else begin
        dirty_29_1 <= _GEN_4242;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_30_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_30_0 <= _GEN_1373;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_30_0 <= _GEN_2302;
      end else begin
        dirty_30_0 <= _GEN_4243;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_30_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_30_1 <= _GEN_1374;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_30_1 <= _GEN_2303;
      end else begin
        dirty_30_1 <= _GEN_4244;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_31_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_31_0 <= _GEN_1375;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_31_0 <= _GEN_2304;
      end else begin
        dirty_31_0 <= _GEN_4245;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_31_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_31_1 <= _GEN_1376;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_31_1 <= _GEN_2305;
      end else begin
        dirty_31_1 <= _GEN_4246;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_32_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_32_0 <= _GEN_1377;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_32_0 <= _GEN_2306;
      end else begin
        dirty_32_0 <= _GEN_4247;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_32_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_32_1 <= _GEN_1378;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_32_1 <= _GEN_2307;
      end else begin
        dirty_32_1 <= _GEN_4248;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_33_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_33_0 <= _GEN_1379;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_33_0 <= _GEN_2308;
      end else begin
        dirty_33_0 <= _GEN_4249;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_33_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_33_1 <= _GEN_1380;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_33_1 <= _GEN_2309;
      end else begin
        dirty_33_1 <= _GEN_4250;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_34_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_34_0 <= _GEN_1381;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_34_0 <= _GEN_2310;
      end else begin
        dirty_34_0 <= _GEN_4251;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_34_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_34_1 <= _GEN_1382;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_34_1 <= _GEN_2311;
      end else begin
        dirty_34_1 <= _GEN_4252;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_35_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_35_0 <= _GEN_1383;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_35_0 <= _GEN_2312;
      end else begin
        dirty_35_0 <= _GEN_4253;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_35_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_35_1 <= _GEN_1384;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_35_1 <= _GEN_2313;
      end else begin
        dirty_35_1 <= _GEN_4254;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_36_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_36_0 <= _GEN_1385;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_36_0 <= _GEN_2314;
      end else begin
        dirty_36_0 <= _GEN_4255;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_36_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_36_1 <= _GEN_1386;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_36_1 <= _GEN_2315;
      end else begin
        dirty_36_1 <= _GEN_4256;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_37_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_37_0 <= _GEN_1387;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_37_0 <= _GEN_2316;
      end else begin
        dirty_37_0 <= _GEN_4257;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_37_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_37_1 <= _GEN_1388;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_37_1 <= _GEN_2317;
      end else begin
        dirty_37_1 <= _GEN_4258;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_38_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_38_0 <= _GEN_1389;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_38_0 <= _GEN_2318;
      end else begin
        dirty_38_0 <= _GEN_4259;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_38_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_38_1 <= _GEN_1390;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_38_1 <= _GEN_2319;
      end else begin
        dirty_38_1 <= _GEN_4260;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_39_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_39_0 <= _GEN_1391;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_39_0 <= _GEN_2320;
      end else begin
        dirty_39_0 <= _GEN_4261;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_39_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_39_1 <= _GEN_1392;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_39_1 <= _GEN_2321;
      end else begin
        dirty_39_1 <= _GEN_4262;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_40_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_40_0 <= _GEN_1393;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_40_0 <= _GEN_2322;
      end else begin
        dirty_40_0 <= _GEN_4263;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_40_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_40_1 <= _GEN_1394;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_40_1 <= _GEN_2323;
      end else begin
        dirty_40_1 <= _GEN_4264;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_41_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_41_0 <= _GEN_1395;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_41_0 <= _GEN_2324;
      end else begin
        dirty_41_0 <= _GEN_4265;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_41_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_41_1 <= _GEN_1396;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_41_1 <= _GEN_2325;
      end else begin
        dirty_41_1 <= _GEN_4266;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_42_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_42_0 <= _GEN_1397;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_42_0 <= _GEN_2326;
      end else begin
        dirty_42_0 <= _GEN_4267;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_42_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_42_1 <= _GEN_1398;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_42_1 <= _GEN_2327;
      end else begin
        dirty_42_1 <= _GEN_4268;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_43_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_43_0 <= _GEN_1399;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_43_0 <= _GEN_2328;
      end else begin
        dirty_43_0 <= _GEN_4269;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_43_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_43_1 <= _GEN_1400;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_43_1 <= _GEN_2329;
      end else begin
        dirty_43_1 <= _GEN_4270;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_44_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_44_0 <= _GEN_1401;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_44_0 <= _GEN_2330;
      end else begin
        dirty_44_0 <= _GEN_4271;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_44_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_44_1 <= _GEN_1402;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_44_1 <= _GEN_2331;
      end else begin
        dirty_44_1 <= _GEN_4272;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_45_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_45_0 <= _GEN_1403;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_45_0 <= _GEN_2332;
      end else begin
        dirty_45_0 <= _GEN_4273;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_45_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_45_1 <= _GEN_1404;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_45_1 <= _GEN_2333;
      end else begin
        dirty_45_1 <= _GEN_4274;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_46_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_46_0 <= _GEN_1405;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_46_0 <= _GEN_2334;
      end else begin
        dirty_46_0 <= _GEN_4275;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_46_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_46_1 <= _GEN_1406;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_46_1 <= _GEN_2335;
      end else begin
        dirty_46_1 <= _GEN_4276;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_47_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_47_0 <= _GEN_1407;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_47_0 <= _GEN_2336;
      end else begin
        dirty_47_0 <= _GEN_4277;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_47_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_47_1 <= _GEN_1408;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_47_1 <= _GEN_2337;
      end else begin
        dirty_47_1 <= _GEN_4278;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_48_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_48_0 <= _GEN_1409;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_48_0 <= _GEN_2338;
      end else begin
        dirty_48_0 <= _GEN_4279;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_48_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_48_1 <= _GEN_1410;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_48_1 <= _GEN_2339;
      end else begin
        dirty_48_1 <= _GEN_4280;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_49_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_49_0 <= _GEN_1411;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_49_0 <= _GEN_2340;
      end else begin
        dirty_49_0 <= _GEN_4281;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_49_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_49_1 <= _GEN_1412;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_49_1 <= _GEN_2341;
      end else begin
        dirty_49_1 <= _GEN_4282;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_50_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_50_0 <= _GEN_1413;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_50_0 <= _GEN_2342;
      end else begin
        dirty_50_0 <= _GEN_4283;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_50_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_50_1 <= _GEN_1414;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_50_1 <= _GEN_2343;
      end else begin
        dirty_50_1 <= _GEN_4284;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_51_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_51_0 <= _GEN_1415;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_51_0 <= _GEN_2344;
      end else begin
        dirty_51_0 <= _GEN_4285;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_51_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_51_1 <= _GEN_1416;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_51_1 <= _GEN_2345;
      end else begin
        dirty_51_1 <= _GEN_4286;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_52_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_52_0 <= _GEN_1417;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_52_0 <= _GEN_2346;
      end else begin
        dirty_52_0 <= _GEN_4287;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_52_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_52_1 <= _GEN_1418;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_52_1 <= _GEN_2347;
      end else begin
        dirty_52_1 <= _GEN_4288;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_53_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_53_0 <= _GEN_1419;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_53_0 <= _GEN_2348;
      end else begin
        dirty_53_0 <= _GEN_4289;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_53_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_53_1 <= _GEN_1420;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_53_1 <= _GEN_2349;
      end else begin
        dirty_53_1 <= _GEN_4290;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_54_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_54_0 <= _GEN_1421;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_54_0 <= _GEN_2350;
      end else begin
        dirty_54_0 <= _GEN_4291;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_54_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_54_1 <= _GEN_1422;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_54_1 <= _GEN_2351;
      end else begin
        dirty_54_1 <= _GEN_4292;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_55_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_55_0 <= _GEN_1423;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_55_0 <= _GEN_2352;
      end else begin
        dirty_55_0 <= _GEN_4293;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_55_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_55_1 <= _GEN_1424;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_55_1 <= _GEN_2353;
      end else begin
        dirty_55_1 <= _GEN_4294;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_56_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_56_0 <= _GEN_1425;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_56_0 <= _GEN_2354;
      end else begin
        dirty_56_0 <= _GEN_4295;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_56_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_56_1 <= _GEN_1426;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_56_1 <= _GEN_2355;
      end else begin
        dirty_56_1 <= _GEN_4296;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_57_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_57_0 <= _GEN_1427;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_57_0 <= _GEN_2356;
      end else begin
        dirty_57_0 <= _GEN_4297;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_57_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_57_1 <= _GEN_1428;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_57_1 <= _GEN_2357;
      end else begin
        dirty_57_1 <= _GEN_4298;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_58_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_58_0 <= _GEN_1429;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_58_0 <= _GEN_2358;
      end else begin
        dirty_58_0 <= _GEN_4299;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_58_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_58_1 <= _GEN_1430;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_58_1 <= _GEN_2359;
      end else begin
        dirty_58_1 <= _GEN_4300;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_59_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_59_0 <= _GEN_1431;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_59_0 <= _GEN_2360;
      end else begin
        dirty_59_0 <= _GEN_4301;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_59_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_59_1 <= _GEN_1432;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_59_1 <= _GEN_2361;
      end else begin
        dirty_59_1 <= _GEN_4302;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_60_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_60_0 <= _GEN_1433;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_60_0 <= _GEN_2362;
      end else begin
        dirty_60_0 <= _GEN_4303;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_60_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_60_1 <= _GEN_1434;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_60_1 <= _GEN_2363;
      end else begin
        dirty_60_1 <= _GEN_4304;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_61_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_61_0 <= _GEN_1435;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_61_0 <= _GEN_2364;
      end else begin
        dirty_61_0 <= _GEN_4305;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_61_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_61_1 <= _GEN_1436;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_61_1 <= _GEN_2365;
      end else begin
        dirty_61_1 <= _GEN_4306;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_62_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_62_0 <= _GEN_1437;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_62_0 <= _GEN_2366;
      end else begin
        dirty_62_0 <= _GEN_4307;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_62_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_62_1 <= _GEN_1438;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_62_1 <= _GEN_2367;
      end else begin
        dirty_62_1 <= _GEN_4308;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_63_0 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_63_0 <= _GEN_1439;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_63_0 <= _GEN_2368;
      end else begin
        dirty_63_0 <= _GEN_4309;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 135:22]
      dirty_63_1 <= 1'h0; // @[playground/src/cache/DCache.scala 135:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          dirty_63_1 <= _GEN_1440;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        dirty_63_1 <= _GEN_2369;
      end else begin
        dirty_63_1 <= _GEN_4310;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_0 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_0 <= _GEN_1249;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_1 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_1 <= _GEN_1250;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_2 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_2 <= _GEN_1251;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_3 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_3 <= _GEN_1252;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_4 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_4 <= _GEN_1253;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_5 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_5 <= _GEN_1254;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_6 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_6 <= _GEN_1255;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_7 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_7 <= _GEN_1256;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_8 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_8 <= _GEN_1257;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_9 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_9 <= _GEN_1258;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_10 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_10 <= _GEN_1259;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_11 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_11 <= _GEN_1260;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_12 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_12 <= _GEN_1261;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_13 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_13 <= _GEN_1262;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_14 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_14 <= _GEN_1263;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_15 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_15 <= _GEN_1264;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_16 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_16 <= _GEN_1265;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_17 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_17 <= _GEN_1266;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_18 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_18 <= _GEN_1267;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_19 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_19 <= _GEN_1268;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_20 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_20 <= _GEN_1269;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_21 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_21 <= _GEN_1270;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_22 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_22 <= _GEN_1271;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_23 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_23 <= _GEN_1272;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_24 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_24 <= _GEN_1273;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_25 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_25 <= _GEN_1274;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_26 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_26 <= _GEN_1275;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_27 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_27 <= _GEN_1276;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_28 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_28 <= _GEN_1277;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_29 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_29 <= _GEN_1278;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_30 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_30 <= _GEN_1279;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_31 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_31 <= _GEN_1280;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_32 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_32 <= _GEN_1281;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_33 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_33 <= _GEN_1282;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_34 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_34 <= _GEN_1283;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_35 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_35 <= _GEN_1284;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_36 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_36 <= _GEN_1285;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_37 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_37 <= _GEN_1286;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_38 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_38 <= _GEN_1287;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_39 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_39 <= _GEN_1288;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_40 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_40 <= _GEN_1289;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_41 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_41 <= _GEN_1290;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_42 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_42 <= _GEN_1291;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_43 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_43 <= _GEN_1292;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_44 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_44 <= _GEN_1293;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_45 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_45 <= _GEN_1294;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_46 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_46 <= _GEN_1295;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_47 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_47 <= _GEN_1296;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_48 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_48 <= _GEN_1297;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_49 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_49 <= _GEN_1298;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_50 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_50 <= _GEN_1299;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_51 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_51 <= _GEN_1300;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_52 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_52 <= _GEN_1301;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_53 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_53 <= _GEN_1302;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_54 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_54 <= _GEN_1303;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_55 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_55 <= _GEN_1304;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_56 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_56 <= _GEN_1305;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_57 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_57 <= _GEN_1306;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_58 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_58 <= _GEN_1307;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_59 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_59 <= _GEN_1308;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_60 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_60 <= _GEN_1309;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_61 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_61 <= _GEN_1310;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_62 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_62 <= _GEN_1311;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 136:22]
      lru_63 <= 1'h0; // @[playground/src/cache/DCache.scala 136:22]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          lru_63 <= _GEN_1312;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 145:22]
      fence <= 1'h0; // @[playground/src/cache/DCache.scala 145:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
          fence <= _GEN_2370;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 148:25]
      readsram <= 1'h0; // @[playground/src/cache/DCache.scala 148:25]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(io_cpu_en)) begin // @[playground/src/cache/DCache.scala 320:23]
        if (io_cpu_fence_i) begin // @[playground/src/cache/DCache.scala 365:30]
          readsram <= _GEN_1650;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
        readsram <= _GEN_2371;
      end else begin
        readsram <= _GEN_4449;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 152:35]
      writeFifo_axi_busy <= 1'h0; // @[playground/src/cache/DCache.scala 152:35]
    end else if (writeFifo_axi_busy) begin // @[playground/src/cache/DCache.scala 290:28]
      if (_T_2) begin // @[playground/src/cache/DCache.scala 298:25]
        writeFifo_axi_busy <= 1'h0; // @[playground/src/cache/DCache.scala 299:26]
      end
    end else begin
      writeFifo_axi_busy <= _GEN_289;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 160:22]
      burst_wstrb_0 <= 8'h0; // @[playground/src/cache/DCache.scala 160:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          burst_wstrb_0 <= _GEN_4315;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 160:22]
      burst_wstrb_1 <= 8'h0; // @[playground/src/cache/DCache.scala 160:22]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          burst_wstrb_1 <= _GEN_4316;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 165:29]
      bank_wbindex <= 3'h0; // @[playground/src/cache/DCache.scala 165:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbindex <= _GEN_2239;
        end else begin
          bank_wbindex <= _GEN_4180;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_0 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_0 <= _GEN_4454;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_1 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_1 <= _GEN_4455;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_2 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_2 <= _GEN_4456;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_3 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_3 <= _GEN_4457;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_4 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_4 <= _GEN_4458;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_5 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_5 <= _GEN_4459;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_6 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_6 <= _GEN_4460;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 166:29]
      bank_wbdata_7 <= 64'h0; // @[playground/src/cache/DCache.scala 166:29]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          bank_wbdata_7 <= _GEN_4461;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 170:30]
      do_replace <= 1'h0; // @[playground/src/cache/DCache.scala 170:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          do_replace <= _GEN_4445;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 567:28]
      ppn <= 20'h0; // @[playground/src/cache/DCache.scala 567:28]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      if (_T_50) begin // @[playground/src/cache/DCache.scala 606:37]
        ppn <= satp_ppn; // @[playground/src/cache/DCache.scala 608:19]
      end
    end else if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
        ppn <= _GEN_5640;
      end else begin
        ppn <= _GEN_5826;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 568:28]
      vpn_index <= 2'h0; // @[playground/src/cache/DCache.scala 568:28]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      if (_T_50) begin // @[playground/src/cache/DCache.scala 606:37]
        vpn_index <= 2'h2; // @[playground/src/cache/DCache.scala 607:19]
      end
    end else if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
        vpn_index <= _GEN_5639;
      end else begin
        vpn_index <= _GEN_5825;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 182:27]
      tag_wstrb_0 <= 1'h0; // @[playground/src/cache/DCache.scala 182:27]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          tag_wstrb_0 <= _GEN_4311;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 182:27]
      tag_wstrb_1 <= 1'h0; // @[playground/src/cache/DCache.scala 182:27]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          tag_wstrb_1 <= _GEN_4312;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 183:27]
      tag_wdata <= 20'h0; // @[playground/src/cache/DCache.scala 183:27]
    end else if (!(3'h0 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
          tag_wdata <= _GEN_4453;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 187:20]
      tag_0 <= 20'h0; // @[playground/src/cache/DCache.scala 187:20]
    end else begin
      tag_0 <= tagRam_0_io_rdata; // @[playground/src/cache/DCache.scala 240:26]
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 187:20]
      tag_1 <= 20'h0; // @[playground/src/cache/DCache.scala 187:20]
    end else begin
      tag_1 <= tagRam_1_io_rdata; // @[playground/src/cache/DCache.scala 240:26]
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 209:28]
      saved_rdata <= 64'h0; // @[playground/src/cache/DCache.scala 209:28]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (io_cpu_en) begin // @[playground/src/cache/DCache.scala 320:23]
        if (!(addr_err)) begin // @[playground/src/cache/DCache.scala 321:24]
          saved_rdata <= _GEN_1441;
        end
      end
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (_T_18) begin // @[playground/src/cache/DCache.scala 383:27]
        saved_rdata <= io_axi_r_bits_data; // @[playground/src/cache/DCache.scala 385:22]
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 259:24]
      ar_addr <= 32'h0; // @[playground/src/cache/DCache.scala 259:24]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      ar_addr <= _GEN_5062;
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      if (pte_uncached) begin // @[playground/src/cache/DCache.scala 622:26]
        ar_addr <= _pte_uncached_T; // @[playground/src/cache/DCache.scala 624:19]
      end else begin
        ar_addr <= _GEN_5062;
      end
    end else begin
      ar_addr <= _GEN_5062;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 259:24]
      ar_len <= 8'h0; // @[playground/src/cache/DCache.scala 259:24]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      ar_len <= _GEN_5063;
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      if (pte_uncached) begin // @[playground/src/cache/DCache.scala 622:26]
        ar_len <= 8'h0; // @[playground/src/cache/DCache.scala 626:19]
      end else begin
        ar_len <= _GEN_5063;
      end
    end else begin
      ar_len <= _GEN_5063;
    end
    ar_size <= _GEN_7927[2:0]; // @[playground/src/cache/DCache.scala 259:{24,24}]
    if (reset) begin // @[playground/src/cache/DCache.scala 260:24]
      arvalid <= 1'h0; // @[playground/src/cache/DCache.scala 260:24]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      arvalid <= _GEN_5065;
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      arvalid <= _GEN_5419;
    end else if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      arvalid <= _GEN_5065;
    end else begin
      arvalid <= _GEN_5809;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 263:23]
      rready <= 1'h0; // @[playground/src/cache/DCache.scala 263:23]
    end else if (3'h0 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      rready <= _GEN_5066;
    end else if (3'h1 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      rready <= _GEN_5423;
    end else if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
      rready <= _GEN_5066;
    end else begin
      rready <= _GEN_5810;
    end
    aw_addr <= _GEN_7928[31:0]; // @[playground/src/cache/DCache.scala 265:{24,24}]
    if (reset) begin // @[playground/src/cache/DCache.scala 265:24]
      aw_len <= 8'h0; // @[playground/src/cache/DCache.scala 265:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      aw_len <= _GEN_299;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      aw_len <= _GEN_299;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      aw_len <= _GEN_2373;
    end else begin
      aw_len <= _GEN_4463;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 265:24]
      aw_size <= 3'h0; // @[playground/src/cache/DCache.scala 265:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      aw_size <= _GEN_296;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      aw_size <= _GEN_296;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      aw_size <= _GEN_2374;
    end else begin
      aw_size <= _GEN_4464;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 266:24]
      awvalid <= 1'h0; // @[playground/src/cache/DCache.scala 266:24]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      awvalid <= _GEN_290;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      awvalid <= _GEN_290;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      awvalid <= _GEN_2237;
    end else begin
      awvalid <= _GEN_4178;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 269:23]
      w_data <= 64'h0; // @[playground/src/cache/DCache.scala 269:23]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_data <= _GEN_297;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_data <= _GEN_297;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_data <= _GEN_2240;
    end else begin
      w_data <= _GEN_4181;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 269:23]
      w_strb <= 8'h0; // @[playground/src/cache/DCache.scala 269:23]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_strb <= _GEN_298;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_strb <= _GEN_298;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_strb <= _GEN_2375;
    end else begin
      w_strb <= _GEN_4465;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 269:23]
      w_last <= 1'h0; // @[playground/src/cache/DCache.scala 269:23]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_last <= _GEN_292;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_last <= _GEN_292;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      w_last <= _GEN_2241;
    end else begin
      w_last <= _GEN_4182;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 270:23]
      wvalid <= 1'h0; // @[playground/src/cache/DCache.scala 270:23]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      wvalid <= _GEN_291;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      wvalid <= _GEN_291;
    end else if (3'h2 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      wvalid <= _GEN_2238;
    end else begin
      wvalid <= _GEN_4179;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 277:29]
      access_fault <= 1'h0; // @[playground/src/cache/DCache.scala 277:29]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      access_fault <= _GEN_1653;
    end else if (3'h1 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      if (_T_18) begin // @[playground/src/cache/DCache.scala 383:27]
        access_fault <= io_axi_r_bits_resp != 2'h0; // @[playground/src/cache/DCache.scala 386:22]
      end
    end else if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      access_fault <= _GEN_4467;
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 278:29]
      page_fault <= 1'h0; // @[playground/src/cache/DCache.scala 278:29]
    end else if (3'h0 == state) begin // @[playground/src/cache/DCache.scala 316:17]
      page_fault <= 1'h0; // @[playground/src/cache/DCache.scala 319:20]
    end else if (!(3'h1 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
      if (!(3'h2 == state)) begin // @[playground/src/cache/DCache.scala 316:17]
        page_fault <= _GEN_4468;
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_ppn <= 20'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_ppn <= _GEN_5629;
        end else begin
          pte_ppn <= _GEN_5815;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_d <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_d <= _GEN_5631;
        end else begin
          pte_flag_d <= _GEN_5817;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_a <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_a <= _GEN_5632;
        end else begin
          pte_flag_a <= _GEN_5818;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_g <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_g <= _GEN_5633;
        end else begin
          pte_flag_g <= _GEN_5819;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_u <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_u <= _GEN_5634;
        end else begin
          pte_flag_u <= _GEN_5820;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_x <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_x <= _GEN_5635;
        end else begin
          pte_flag_x <= _GEN_5821;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_w <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_w <= _GEN_5636;
        end else begin
          pte_flag_w <= _GEN_5822;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_r <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_r <= _GEN_5637;
        end else begin
          pte_flag_r <= _GEN_5823;
        end
      end
    end
    if (reset) begin // @[playground/src/cache/DCache.scala 569:28]
      pte_flag_v <= 1'h0; // @[playground/src/cache/DCache.scala 569:28]
    end else if (!(3'h0 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
      if (!(3'h1 == ptw_state)) begin // @[playground/src/cache/DCache.scala 603:21]
        if (3'h2 == ptw_state) begin // @[playground/src/cache/DCache.scala 603:21]
          pte_flag_v <= _GEN_5638;
        end else begin
          pte_flag_v <= _GEN_5824;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ptw_state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  ptw_scratch_paddr_tag = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  ptw_scratch_paddr_index = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  ptw_scratch_paddr_offset = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  ptw_scratch_replace = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ptw_scratch_dcache_wait = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_0_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_0_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_1_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_1_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_2_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_2_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_3_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_3_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_4_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_4_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_5_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_5_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_6_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_6_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_7_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_7_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_8_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_8_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_9_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_9_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_10_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_10_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_11_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_11_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_12_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_12_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_13_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_13_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_14_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_14_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_15_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_15_1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_16_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_16_1 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_17_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_17_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_18_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_18_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_19_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_19_1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_20_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_20_1 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_21_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_21_1 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_22_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_22_1 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_23_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_23_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_24_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_24_1 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_25_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_25_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_26_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_26_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_27_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_27_1 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_28_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_28_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_29_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_29_1 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_30_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_30_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_31_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_31_1 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_32_0 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_32_1 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_33_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_33_1 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_34_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_34_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_35_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_35_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_36_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_36_1 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_37_0 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_37_1 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_38_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_38_1 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_39_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_39_1 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_40_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_40_1 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_41_0 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_41_1 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_42_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_42_1 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_43_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_43_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_44_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_44_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_45_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_45_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_46_0 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_46_1 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_47_0 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_47_1 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_48_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_48_1 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_49_0 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_49_1 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_50_0 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_50_1 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_51_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_51_1 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_52_0 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_52_1 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_53_0 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_53_1 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_54_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_54_1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_55_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_55_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_56_0 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_56_1 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_57_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_57_1 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_58_0 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_58_1 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_59_0 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_59_1 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_60_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_60_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_61_0 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_61_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_62_0 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_62_1 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_63_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_63_1 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  dirty_0_0 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  dirty_0_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dirty_1_0 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  dirty_1_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  dirty_2_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dirty_2_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  dirty_3_0 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  dirty_3_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dirty_4_0 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  dirty_4_1 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  dirty_5_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dirty_5_1 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  dirty_6_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  dirty_6_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dirty_7_0 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  dirty_7_1 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  dirty_8_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dirty_8_1 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  dirty_9_0 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dirty_9_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dirty_10_0 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dirty_10_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  dirty_11_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dirty_11_1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  dirty_12_0 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dirty_12_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dirty_13_0 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dirty_13_1 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  dirty_14_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dirty_14_1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  dirty_15_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dirty_15_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dirty_16_0 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dirty_16_1 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  dirty_17_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dirty_17_1 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  dirty_18_0 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dirty_18_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dirty_19_0 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dirty_19_1 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  dirty_20_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dirty_20_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  dirty_21_0 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dirty_21_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dirty_22_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dirty_22_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  dirty_23_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dirty_23_1 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  dirty_24_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dirty_24_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dirty_25_0 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  dirty_25_1 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  dirty_26_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dirty_26_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  dirty_27_0 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  dirty_27_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dirty_28_0 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_28_1 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_29_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_29_1 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_30_0 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dirty_30_1 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dirty_31_0 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dirty_31_1 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dirty_32_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dirty_32_1 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dirty_33_0 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dirty_33_1 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dirty_34_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dirty_34_1 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dirty_35_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dirty_35_1 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dirty_36_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dirty_36_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dirty_37_0 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dirty_37_1 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dirty_38_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dirty_38_1 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dirty_39_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dirty_39_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dirty_40_0 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dirty_40_1 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  dirty_41_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dirty_41_1 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  dirty_42_0 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dirty_42_1 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dirty_43_0 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dirty_43_1 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  dirty_44_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dirty_44_1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  dirty_45_0 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  dirty_45_1 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dirty_46_0 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  dirty_46_1 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  dirty_47_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dirty_47_1 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  dirty_48_0 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  dirty_48_1 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dirty_49_0 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  dirty_49_1 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  dirty_50_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dirty_50_1 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  dirty_51_0 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  dirty_51_1 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dirty_52_0 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  dirty_52_1 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  dirty_53_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dirty_53_1 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  dirty_54_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  dirty_54_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dirty_55_0 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  dirty_55_1 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  dirty_56_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dirty_56_1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  dirty_57_0 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  dirty_57_1 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dirty_58_0 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dirty_58_1 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  dirty_59_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dirty_59_1 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  dirty_60_0 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  dirty_60_1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  dirty_61_0 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  dirty_61_1 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  dirty_62_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dirty_62_1 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  dirty_63_0 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  dirty_63_1 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  lru_0 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  lru_1 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  lru_2 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  lru_3 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  lru_4 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  lru_5 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  lru_6 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  lru_7 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  lru_8 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  lru_9 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  lru_10 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  lru_11 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  lru_12 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  lru_13 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  lru_14 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  lru_15 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  lru_16 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  lru_17 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  lru_18 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  lru_19 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  lru_20 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  lru_21 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  lru_22 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  lru_23 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  lru_24 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  lru_25 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  lru_26 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  lru_27 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  lru_28 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  lru_29 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  lru_30 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  lru_31 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  lru_32 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  lru_33 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  lru_34 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  lru_35 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  lru_36 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  lru_37 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  lru_38 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  lru_39 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  lru_40 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  lru_41 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  lru_42 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  lru_43 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  lru_44 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  lru_45 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  lru_46 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  lru_47 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  lru_48 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  lru_49 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  lru_50 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  lru_51 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  lru_52 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  lru_53 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  lru_54 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  lru_55 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  lru_56 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  lru_57 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  lru_58 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  lru_59 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  lru_60 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  lru_61 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  lru_62 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  lru_63 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  fence = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  readsram = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  writeFifo_axi_busy = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  burst_wstrb_0 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  burst_wstrb_1 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  bank_wbindex = _RAND_332[2:0];
  _RAND_333 = {2{`RANDOM}};
  bank_wbdata_0 = _RAND_333[63:0];
  _RAND_334 = {2{`RANDOM}};
  bank_wbdata_1 = _RAND_334[63:0];
  _RAND_335 = {2{`RANDOM}};
  bank_wbdata_2 = _RAND_335[63:0];
  _RAND_336 = {2{`RANDOM}};
  bank_wbdata_3 = _RAND_336[63:0];
  _RAND_337 = {2{`RANDOM}};
  bank_wbdata_4 = _RAND_337[63:0];
  _RAND_338 = {2{`RANDOM}};
  bank_wbdata_5 = _RAND_338[63:0];
  _RAND_339 = {2{`RANDOM}};
  bank_wbdata_6 = _RAND_339[63:0];
  _RAND_340 = {2{`RANDOM}};
  bank_wbdata_7 = _RAND_340[63:0];
  _RAND_341 = {1{`RANDOM}};
  do_replace = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ppn = _RAND_342[19:0];
  _RAND_343 = {1{`RANDOM}};
  vpn_index = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  tag_wstrb_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  tag_wstrb_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  tag_wdata = _RAND_346[19:0];
  _RAND_347 = {1{`RANDOM}};
  tag_0 = _RAND_347[19:0];
  _RAND_348 = {1{`RANDOM}};
  tag_1 = _RAND_348[19:0];
  _RAND_349 = {2{`RANDOM}};
  saved_rdata = _RAND_349[63:0];
  _RAND_350 = {1{`RANDOM}};
  ar_addr = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  ar_len = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  ar_size = _RAND_352[2:0];
  _RAND_353 = {1{`RANDOM}};
  arvalid = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  rready = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  aw_addr = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  aw_len = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  aw_size = _RAND_357[2:0];
  _RAND_358 = {1{`RANDOM}};
  awvalid = _RAND_358[0:0];
  _RAND_359 = {2{`RANDOM}};
  w_data = _RAND_359[63:0];
  _RAND_360 = {1{`RANDOM}};
  w_strb = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  w_last = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  wvalid = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  access_fault = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  page_fault = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  pte_ppn = _RAND_365[19:0];
  _RAND_366 = {1{`RANDOM}};
  pte_flag_d = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  pte_flag_a = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  pte_flag_g = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  pte_flag_u = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  pte_flag_x = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  pte_flag_w = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  pte_flag_r = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  pte_flag_v = _RAND_373[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheAXIInterface(
  input         clock,
  input         reset,
  output        io_icache_ar_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_icache_ar_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [31:0] io_icache_ar_bits_addr, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [7:0]  io_icache_ar_bits_len, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [2:0]  io_icache_ar_bits_size, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_icache_r_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_icache_r_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [63:0] io_icache_r_bits_data, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [1:0]  io_icache_r_bits_resp, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_icache_r_bits_last, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_dcache_ar_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_dcache_ar_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [31:0] io_dcache_ar_bits_addr, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [7:0]  io_dcache_ar_bits_len, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [2:0]  io_dcache_ar_bits_size, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_dcache_r_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_dcache_r_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [63:0] io_dcache_r_bits_data, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [1:0]  io_dcache_r_bits_resp, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_dcache_r_bits_last, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_dcache_aw_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_dcache_aw_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [31:0] io_dcache_aw_bits_addr, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [7:0]  io_dcache_aw_bits_len, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [2:0]  io_dcache_aw_bits_size, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_dcache_w_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_dcache_w_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [63:0] io_dcache_w_bits_data, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [7:0]  io_dcache_w_bits_strb, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_dcache_w_bits_last, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_dcache_b_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_axi_ar_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_axi_ar_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [3:0]  io_axi_ar_bits_id, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [31:0] io_axi_ar_bits_addr, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [7:0]  io_axi_ar_bits_len, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [2:0]  io_axi_ar_bits_size, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_axi_r_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_axi_r_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [3:0]  io_axi_r_bits_id, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [63:0] io_axi_r_bits_data, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input  [1:0]  io_axi_r_bits_resp, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_axi_r_bits_last, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_axi_aw_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_axi_aw_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [31:0] io_axi_aw_bits_addr, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [7:0]  io_axi_aw_bits_len, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [2:0]  io_axi_aw_bits_size, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_axi_w_ready, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_axi_w_valid, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [63:0] io_axi_w_bits_data, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output [7:0]  io_axi_w_bits_strb, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  output        io_axi_w_bits_last, // @[playground/src/cache/CacheAXIInterface.scala 8:14]
  input         io_axi_b_valid // @[playground/src/cache/CacheAXIInterface.scala 8:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  ar_sel_lock; // @[playground/src/cache/CacheAXIInterface.scala 45:30]
  reg  ar_sel_val; // @[playground/src/cache/CacheAXIInterface.scala 46:30]
  wire  choose_dcache = ar_sel_lock ? ar_sel_val : ~io_icache_ar_valid & io_dcache_ar_valid; // @[playground/src/cache/CacheAXIInterface.scala 47:26]
  wire  r_sel = io_axi_r_bits_id[0]; // @[playground/src/cache/CacheAXIInterface.scala 72:31]
  assign io_icache_ar_ready = ~choose_dcache & io_axi_ar_ready; // @[playground/src/cache/CacheAXIInterface.scala 67:42]
  assign io_icache_r_valid = ~r_sel & io_axi_r_valid; // @[playground/src/cache/CacheAXIInterface.scala 77:35]
  assign io_icache_r_bits_data = io_axi_r_bits_data; // @[playground/src/cache/CacheAXIInterface.scala 74:25]
  assign io_icache_r_bits_resp = io_axi_r_bits_resp; // @[playground/src/cache/CacheAXIInterface.scala 75:25]
  assign io_icache_r_bits_last = io_axi_r_bits_last; // @[playground/src/cache/CacheAXIInterface.scala 76:25]
  assign io_dcache_ar_ready = choose_dcache & io_axi_ar_ready; // @[playground/src/cache/CacheAXIInterface.scala 68:41]
  assign io_dcache_r_valid = r_sel & io_axi_r_valid; // @[playground/src/cache/CacheAXIInterface.scala 82:34]
  assign io_dcache_r_bits_data = io_axi_r_bits_data; // @[playground/src/cache/CacheAXIInterface.scala 79:25]
  assign io_dcache_r_bits_resp = io_axi_r_bits_resp; // @[playground/src/cache/CacheAXIInterface.scala 80:25]
  assign io_dcache_r_bits_last = io_axi_r_bits_last; // @[playground/src/cache/CacheAXIInterface.scala 81:25]
  assign io_dcache_aw_ready = io_axi_aw_ready; // @[playground/src/cache/CacheAXIInterface.scala 24:24]
  assign io_dcache_w_ready = io_axi_w_ready; // @[playground/src/cache/CacheAXIInterface.scala 33:22]
  assign io_dcache_b_valid = io_axi_b_valid; // @[playground/src/cache/CacheAXIInterface.scala 38:25]
  assign io_axi_ar_valid = choose_dcache ? io_dcache_ar_valid : io_icache_ar_valid; // @[playground/src/cache/CacheAXIInterface.scala 62:30]
  assign io_axi_ar_bits_id = {3'h0,choose_dcache}; // @[playground/src/cache/CacheAXIInterface.scala 58:30]
  assign io_axi_ar_bits_addr = choose_dcache ? io_dcache_ar_bits_addr : io_icache_ar_bits_addr; // @[playground/src/cache/CacheAXIInterface.scala 59:30]
  assign io_axi_ar_bits_len = choose_dcache ? io_dcache_ar_bits_len : io_icache_ar_bits_len; // @[playground/src/cache/CacheAXIInterface.scala 60:30]
  assign io_axi_ar_bits_size = choose_dcache ? io_dcache_ar_bits_size : io_icache_ar_bits_size; // @[playground/src/cache/CacheAXIInterface.scala 61:30]
  assign io_axi_r_ready = r_sel ? io_dcache_r_ready : io_icache_r_ready; // @[playground/src/cache/CacheAXIInterface.scala 83:31]
  assign io_axi_aw_valid = io_dcache_aw_valid; // @[playground/src/cache/CacheAXIInterface.scala 19:24]
  assign io_axi_aw_bits_addr = io_dcache_aw_bits_addr; // @[playground/src/cache/CacheAXIInterface.scala 16:24]
  assign io_axi_aw_bits_len = io_dcache_aw_bits_len; // @[playground/src/cache/CacheAXIInterface.scala 17:24]
  assign io_axi_aw_bits_size = io_dcache_aw_bits_size; // @[playground/src/cache/CacheAXIInterface.scala 18:24]
  assign io_axi_w_valid = io_dcache_w_valid; // @[playground/src/cache/CacheAXIInterface.scala 32:22]
  assign io_axi_w_bits_data = io_dcache_w_bits_data; // @[playground/src/cache/CacheAXIInterface.scala 29:22]
  assign io_axi_w_bits_strb = io_dcache_w_bits_strb; // @[playground/src/cache/CacheAXIInterface.scala 30:22]
  assign io_axi_w_bits_last = io_dcache_w_bits_last; // @[playground/src/cache/CacheAXIInterface.scala 31:22]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/cache/CacheAXIInterface.scala 45:30]
      ar_sel_lock <= 1'h0; // @[playground/src/cache/CacheAXIInterface.scala 45:30]
    end else if (io_axi_ar_valid) begin // @[playground/src/cache/CacheAXIInterface.scala 49:25]
      if (io_axi_ar_ready) begin // @[playground/src/cache/CacheAXIInterface.scala 50:27]
        ar_sel_lock <= 1'h0; // @[playground/src/cache/CacheAXIInterface.scala 51:19]
      end else begin
        ar_sel_lock <= 1'h1; // @[playground/src/cache/CacheAXIInterface.scala 53:19]
      end
    end
    if (reset) begin // @[playground/src/cache/CacheAXIInterface.scala 46:30]
      ar_sel_val <= 1'h0; // @[playground/src/cache/CacheAXIInterface.scala 46:30]
    end else if (io_axi_ar_valid) begin // @[playground/src/cache/CacheAXIInterface.scala 49:25]
      if (!(io_axi_ar_ready)) begin // @[playground/src/cache/CacheAXIInterface.scala 50:27]
        if (!(ar_sel_lock)) begin // @[playground/src/cache/CacheAXIInterface.scala 47:26]
          ar_sel_val <= ~io_icache_ar_valid & io_dcache_ar_valid;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_sel_lock = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ar_sel_val = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache(
  input         clock,
  input         reset,
  input         io_inst_req, // @[playground/src/cache/Cache.scala 11:14]
  input         io_inst_complete_single_request, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_inst_addr_0, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_inst_addr_1, // @[playground/src/cache/Cache.scala 11:14]
  input         io_inst_fence_i, // @[playground/src/cache/Cache.scala 11:14]
  input         io_inst_dcache_stall, // @[playground/src/cache/Cache.scala 11:14]
  output [63:0] io_inst_inst_0, // @[playground/src/cache/Cache.scala 11:14]
  output [63:0] io_inst_inst_1, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_inst_valid_0, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_inst_valid_1, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_access_fault, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_page_fault, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_addr_misaligned, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_icache_stall, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_tlb_en, // @[playground/src/cache/Cache.scala 11:14]
  output [63:0] io_inst_tlb_vaddr, // @[playground/src/cache/Cache.scala 11:14]
  output        io_inst_tlb_complete_single_request, // @[playground/src/cache/Cache.scala 11:14]
  input         io_inst_tlb_uncached, // @[playground/src/cache/Cache.scala 11:14]
  input         io_inst_tlb_hit, // @[playground/src/cache/Cache.scala 11:14]
  input  [19:0] io_inst_tlb_ptag, // @[playground/src/cache/Cache.scala 11:14]
  input  [31:0] io_inst_tlb_paddr, // @[playground/src/cache/Cache.scala 11:14]
  input         io_inst_tlb_page_fault, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_data_exe_addr, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_data_addr, // @[playground/src/cache/Cache.scala 11:14]
  input  [7:0]  io_data_rlen, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_en, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_wen, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_data_wdata, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_complete_single_request, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_fence_i, // @[playground/src/cache/Cache.scala 11:14]
  input  [7:0]  io_data_wstrb, // @[playground/src/cache/Cache.scala 11:14]
  output [63:0] io_data_rdata, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_access_fault, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_page_fault, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_dcache_ready, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_en, // @[playground/src/cache/Cache.scala 11:14]
  output [63:0] io_data_tlb_vaddr, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_complete_single_request, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_tlb_uncached, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_tlb_hit, // @[playground/src/cache/Cache.scala 11:14]
  input  [19:0] io_data_tlb_ptag, // @[playground/src/cache/Cache.scala 11:14]
  input  [31:0] io_data_tlb_paddr, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_tlb_page_fault, // @[playground/src/cache/Cache.scala 11:14]
  output [1:0]  io_data_tlb_access_type, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_vpn_ready, // @[playground/src/cache/Cache.scala 11:14]
  input         io_data_tlb_ptw_vpn_valid, // @[playground/src/cache/Cache.scala 11:14]
  input  [26:0] io_data_tlb_ptw_vpn_bits, // @[playground/src/cache/Cache.scala 11:14]
  input  [1:0]  io_data_tlb_ptw_access_type, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_valid, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_page_fault, // @[playground/src/cache/Cache.scala 11:14]
  output [19:0] io_data_tlb_ptw_pte_bits_entry_ppn, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_d, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_g, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_u, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_x, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_w, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_r, // @[playground/src/cache/Cache.scala 11:14]
  output        io_data_tlb_ptw_pte_bits_entry_flag_v, // @[playground/src/cache/Cache.scala 11:14]
  output [17:0] io_data_tlb_ptw_pte_bits_rmask, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_data_tlb_csr_satp, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_data_tlb_csr_mstatus, // @[playground/src/cache/Cache.scala 11:14]
  input  [1:0]  io_data_tlb_csr_imode, // @[playground/src/cache/Cache.scala 11:14]
  input  [1:0]  io_data_tlb_csr_dmode, // @[playground/src/cache/Cache.scala 11:14]
  input         io_axi_ar_ready, // @[playground/src/cache/Cache.scala 11:14]
  output        io_axi_ar_valid, // @[playground/src/cache/Cache.scala 11:14]
  output [3:0]  io_axi_ar_bits_id, // @[playground/src/cache/Cache.scala 11:14]
  output [31:0] io_axi_ar_bits_addr, // @[playground/src/cache/Cache.scala 11:14]
  output [7:0]  io_axi_ar_bits_len, // @[playground/src/cache/Cache.scala 11:14]
  output [2:0]  io_axi_ar_bits_size, // @[playground/src/cache/Cache.scala 11:14]
  output        io_axi_r_ready, // @[playground/src/cache/Cache.scala 11:14]
  input         io_axi_r_valid, // @[playground/src/cache/Cache.scala 11:14]
  input  [3:0]  io_axi_r_bits_id, // @[playground/src/cache/Cache.scala 11:14]
  input  [63:0] io_axi_r_bits_data, // @[playground/src/cache/Cache.scala 11:14]
  input  [1:0]  io_axi_r_bits_resp, // @[playground/src/cache/Cache.scala 11:14]
  input         io_axi_r_bits_last, // @[playground/src/cache/Cache.scala 11:14]
  input         io_axi_aw_ready, // @[playground/src/cache/Cache.scala 11:14]
  output        io_axi_aw_valid, // @[playground/src/cache/Cache.scala 11:14]
  output [31:0] io_axi_aw_bits_addr, // @[playground/src/cache/Cache.scala 11:14]
  output [7:0]  io_axi_aw_bits_len, // @[playground/src/cache/Cache.scala 11:14]
  output [2:0]  io_axi_aw_bits_size, // @[playground/src/cache/Cache.scala 11:14]
  input         io_axi_w_ready, // @[playground/src/cache/Cache.scala 11:14]
  output        io_axi_w_valid, // @[playground/src/cache/Cache.scala 11:14]
  output [63:0] io_axi_w_bits_data, // @[playground/src/cache/Cache.scala 11:14]
  output [7:0]  io_axi_w_bits_strb, // @[playground/src/cache/Cache.scala 11:14]
  output        io_axi_w_bits_last, // @[playground/src/cache/Cache.scala 11:14]
  input         io_axi_b_valid // @[playground/src/cache/Cache.scala 11:14]
);
  wire  icache_clock; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_reset; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_req; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_complete_single_request; // @[playground/src/cache/Cache.scala 20:29]
  wire [63:0] icache_io_cpu_addr_0; // @[playground/src/cache/Cache.scala 20:29]
  wire [63:0] icache_io_cpu_addr_1; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_fence_i; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_dcache_stall; // @[playground/src/cache/Cache.scala 20:29]
  wire [63:0] icache_io_cpu_inst_0; // @[playground/src/cache/Cache.scala 20:29]
  wire [63:0] icache_io_cpu_inst_1; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_inst_valid_0; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_inst_valid_1; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_access_fault; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_page_fault; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_addr_misaligned; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_icache_stall; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_tlb_en; // @[playground/src/cache/Cache.scala 20:29]
  wire [63:0] icache_io_cpu_tlb_vaddr; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_tlb_complete_single_request; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_tlb_uncached; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_tlb_hit; // @[playground/src/cache/Cache.scala 20:29]
  wire [19:0] icache_io_cpu_tlb_ptag; // @[playground/src/cache/Cache.scala 20:29]
  wire [31:0] icache_io_cpu_tlb_paddr; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_cpu_tlb_page_fault; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_axi_ar_ready; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_axi_ar_valid; // @[playground/src/cache/Cache.scala 20:29]
  wire [31:0] icache_io_axi_ar_bits_addr; // @[playground/src/cache/Cache.scala 20:29]
  wire [7:0] icache_io_axi_ar_bits_len; // @[playground/src/cache/Cache.scala 20:29]
  wire [2:0] icache_io_axi_ar_bits_size; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_axi_r_ready; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_axi_r_valid; // @[playground/src/cache/Cache.scala 20:29]
  wire [63:0] icache_io_axi_r_bits_data; // @[playground/src/cache/Cache.scala 20:29]
  wire [1:0] icache_io_axi_r_bits_resp; // @[playground/src/cache/Cache.scala 20:29]
  wire  icache_io_axi_r_bits_last; // @[playground/src/cache/Cache.scala 20:29]
  wire  dcache_clock; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_reset; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_exe_addr; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_addr; // @[playground/src/cache/Cache.scala 21:29]
  wire [7:0] dcache_io_cpu_rlen; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_en; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_wen; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_wdata; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_complete_single_request; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_fence_i; // @[playground/src/cache/Cache.scala 21:29]
  wire [7:0] dcache_io_cpu_wstrb; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_rdata; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_access_fault; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_page_fault; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_dcache_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_en; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_tlb_vaddr; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_complete_single_request; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_uncached; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_hit; // @[playground/src/cache/Cache.scala 21:29]
  wire [19:0] dcache_io_cpu_tlb_ptag; // @[playground/src/cache/Cache.scala 21:29]
  wire [31:0] dcache_io_cpu_tlb_paddr; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_page_fault; // @[playground/src/cache/Cache.scala 21:29]
  wire [1:0] dcache_io_cpu_tlb_access_type; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_vpn_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_vpn_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire [26:0] dcache_io_cpu_tlb_ptw_vpn_bits; // @[playground/src/cache/Cache.scala 21:29]
  wire [1:0] dcache_io_cpu_tlb_ptw_access_type; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_access_fault; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_page_fault; // @[playground/src/cache/Cache.scala 21:29]
  wire [19:0] dcache_io_cpu_tlb_ptw_pte_bits_entry_ppn; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_d; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_g; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_u; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_x; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_w; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_r; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_v; // @[playground/src/cache/Cache.scala 21:29]
  wire [17:0] dcache_io_cpu_tlb_ptw_pte_bits_rmask; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_tlb_csr_satp; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_cpu_tlb_csr_mstatus; // @[playground/src/cache/Cache.scala 21:29]
  wire [1:0] dcache_io_cpu_tlb_csr_imode; // @[playground/src/cache/Cache.scala 21:29]
  wire [1:0] dcache_io_cpu_tlb_csr_dmode; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_ar_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_ar_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire [31:0] dcache_io_axi_ar_bits_addr; // @[playground/src/cache/Cache.scala 21:29]
  wire [7:0] dcache_io_axi_ar_bits_len; // @[playground/src/cache/Cache.scala 21:29]
  wire [2:0] dcache_io_axi_ar_bits_size; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_r_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_r_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_axi_r_bits_data; // @[playground/src/cache/Cache.scala 21:29]
  wire [1:0] dcache_io_axi_r_bits_resp; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_r_bits_last; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_aw_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_aw_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire [31:0] dcache_io_axi_aw_bits_addr; // @[playground/src/cache/Cache.scala 21:29]
  wire [7:0] dcache_io_axi_aw_bits_len; // @[playground/src/cache/Cache.scala 21:29]
  wire [2:0] dcache_io_axi_aw_bits_size; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_w_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_w_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire [63:0] dcache_io_axi_w_bits_data; // @[playground/src/cache/Cache.scala 21:29]
  wire [7:0] dcache_io_axi_w_bits_strb; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_w_bits_last; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_b_ready; // @[playground/src/cache/Cache.scala 21:29]
  wire  dcache_io_axi_b_valid; // @[playground/src/cache/Cache.scala 21:29]
  wire  axi_interface_clock; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_reset; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_icache_ar_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_icache_ar_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [31:0] axi_interface_io_icache_ar_bits_addr; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_icache_ar_bits_len; // @[playground/src/cache/Cache.scala 22:29]
  wire [2:0] axi_interface_io_icache_ar_bits_size; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_icache_r_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_icache_r_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [63:0] axi_interface_io_icache_r_bits_data; // @[playground/src/cache/Cache.scala 22:29]
  wire [1:0] axi_interface_io_icache_r_bits_resp; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_icache_r_bits_last; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_ar_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_ar_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [31:0] axi_interface_io_dcache_ar_bits_addr; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_dcache_ar_bits_len; // @[playground/src/cache/Cache.scala 22:29]
  wire [2:0] axi_interface_io_dcache_ar_bits_size; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_r_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_r_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [63:0] axi_interface_io_dcache_r_bits_data; // @[playground/src/cache/Cache.scala 22:29]
  wire [1:0] axi_interface_io_dcache_r_bits_resp; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_r_bits_last; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_aw_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_aw_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [31:0] axi_interface_io_dcache_aw_bits_addr; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_dcache_aw_bits_len; // @[playground/src/cache/Cache.scala 22:29]
  wire [2:0] axi_interface_io_dcache_aw_bits_size; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_w_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_w_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [63:0] axi_interface_io_dcache_w_bits_data; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_dcache_w_bits_strb; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_w_bits_last; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_dcache_b_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_ar_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_ar_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [3:0] axi_interface_io_axi_ar_bits_id; // @[playground/src/cache/Cache.scala 22:29]
  wire [31:0] axi_interface_io_axi_ar_bits_addr; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_axi_ar_bits_len; // @[playground/src/cache/Cache.scala 22:29]
  wire [2:0] axi_interface_io_axi_ar_bits_size; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_r_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_r_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [3:0] axi_interface_io_axi_r_bits_id; // @[playground/src/cache/Cache.scala 22:29]
  wire [63:0] axi_interface_io_axi_r_bits_data; // @[playground/src/cache/Cache.scala 22:29]
  wire [1:0] axi_interface_io_axi_r_bits_resp; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_r_bits_last; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_aw_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_aw_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [31:0] axi_interface_io_axi_aw_bits_addr; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_axi_aw_bits_len; // @[playground/src/cache/Cache.scala 22:29]
  wire [2:0] axi_interface_io_axi_aw_bits_size; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_w_ready; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_w_valid; // @[playground/src/cache/Cache.scala 22:29]
  wire [63:0] axi_interface_io_axi_w_bits_data; // @[playground/src/cache/Cache.scala 22:29]
  wire [7:0] axi_interface_io_axi_w_bits_strb; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_w_bits_last; // @[playground/src/cache/Cache.scala 22:29]
  wire  axi_interface_io_axi_b_valid; // @[playground/src/cache/Cache.scala 22:29]
  ICache icache ( // @[playground/src/cache/Cache.scala 20:29]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_cpu_req(icache_io_cpu_req),
    .io_cpu_complete_single_request(icache_io_cpu_complete_single_request),
    .io_cpu_addr_0(icache_io_cpu_addr_0),
    .io_cpu_addr_1(icache_io_cpu_addr_1),
    .io_cpu_fence_i(icache_io_cpu_fence_i),
    .io_cpu_dcache_stall(icache_io_cpu_dcache_stall),
    .io_cpu_inst_0(icache_io_cpu_inst_0),
    .io_cpu_inst_1(icache_io_cpu_inst_1),
    .io_cpu_inst_valid_0(icache_io_cpu_inst_valid_0),
    .io_cpu_inst_valid_1(icache_io_cpu_inst_valid_1),
    .io_cpu_access_fault(icache_io_cpu_access_fault),
    .io_cpu_page_fault(icache_io_cpu_page_fault),
    .io_cpu_addr_misaligned(icache_io_cpu_addr_misaligned),
    .io_cpu_icache_stall(icache_io_cpu_icache_stall),
    .io_cpu_tlb_en(icache_io_cpu_tlb_en),
    .io_cpu_tlb_vaddr(icache_io_cpu_tlb_vaddr),
    .io_cpu_tlb_complete_single_request(icache_io_cpu_tlb_complete_single_request),
    .io_cpu_tlb_uncached(icache_io_cpu_tlb_uncached),
    .io_cpu_tlb_hit(icache_io_cpu_tlb_hit),
    .io_cpu_tlb_ptag(icache_io_cpu_tlb_ptag),
    .io_cpu_tlb_paddr(icache_io_cpu_tlb_paddr),
    .io_cpu_tlb_page_fault(icache_io_cpu_tlb_page_fault),
    .io_axi_ar_ready(icache_io_axi_ar_ready),
    .io_axi_ar_valid(icache_io_axi_ar_valid),
    .io_axi_ar_bits_addr(icache_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(icache_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(icache_io_axi_ar_bits_size),
    .io_axi_r_ready(icache_io_axi_r_ready),
    .io_axi_r_valid(icache_io_axi_r_valid),
    .io_axi_r_bits_data(icache_io_axi_r_bits_data),
    .io_axi_r_bits_resp(icache_io_axi_r_bits_resp),
    .io_axi_r_bits_last(icache_io_axi_r_bits_last)
  );
  DCache dcache ( // @[playground/src/cache/Cache.scala 21:29]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_cpu_exe_addr(dcache_io_cpu_exe_addr),
    .io_cpu_addr(dcache_io_cpu_addr),
    .io_cpu_rlen(dcache_io_cpu_rlen),
    .io_cpu_en(dcache_io_cpu_en),
    .io_cpu_wen(dcache_io_cpu_wen),
    .io_cpu_wdata(dcache_io_cpu_wdata),
    .io_cpu_complete_single_request(dcache_io_cpu_complete_single_request),
    .io_cpu_fence_i(dcache_io_cpu_fence_i),
    .io_cpu_wstrb(dcache_io_cpu_wstrb),
    .io_cpu_rdata(dcache_io_cpu_rdata),
    .io_cpu_access_fault(dcache_io_cpu_access_fault),
    .io_cpu_page_fault(dcache_io_cpu_page_fault),
    .io_cpu_dcache_ready(dcache_io_cpu_dcache_ready),
    .io_cpu_tlb_en(dcache_io_cpu_tlb_en),
    .io_cpu_tlb_vaddr(dcache_io_cpu_tlb_vaddr),
    .io_cpu_tlb_complete_single_request(dcache_io_cpu_tlb_complete_single_request),
    .io_cpu_tlb_uncached(dcache_io_cpu_tlb_uncached),
    .io_cpu_tlb_hit(dcache_io_cpu_tlb_hit),
    .io_cpu_tlb_ptag(dcache_io_cpu_tlb_ptag),
    .io_cpu_tlb_paddr(dcache_io_cpu_tlb_paddr),
    .io_cpu_tlb_page_fault(dcache_io_cpu_tlb_page_fault),
    .io_cpu_tlb_access_type(dcache_io_cpu_tlb_access_type),
    .io_cpu_tlb_ptw_vpn_ready(dcache_io_cpu_tlb_ptw_vpn_ready),
    .io_cpu_tlb_ptw_vpn_valid(dcache_io_cpu_tlb_ptw_vpn_valid),
    .io_cpu_tlb_ptw_vpn_bits(dcache_io_cpu_tlb_ptw_vpn_bits),
    .io_cpu_tlb_ptw_access_type(dcache_io_cpu_tlb_ptw_access_type),
    .io_cpu_tlb_ptw_pte_valid(dcache_io_cpu_tlb_ptw_pte_valid),
    .io_cpu_tlb_ptw_pte_bits_access_fault(dcache_io_cpu_tlb_ptw_pte_bits_access_fault),
    .io_cpu_tlb_ptw_pte_bits_page_fault(dcache_io_cpu_tlb_ptw_pte_bits_page_fault),
    .io_cpu_tlb_ptw_pte_bits_entry_ppn(dcache_io_cpu_tlb_ptw_pte_bits_entry_ppn),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_d(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_d),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_g(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_g),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_u(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_u),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_x(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_x),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_w(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_w),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_r(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_r),
    .io_cpu_tlb_ptw_pte_bits_entry_flag_v(dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_v),
    .io_cpu_tlb_ptw_pte_bits_rmask(dcache_io_cpu_tlb_ptw_pte_bits_rmask),
    .io_cpu_tlb_csr_satp(dcache_io_cpu_tlb_csr_satp),
    .io_cpu_tlb_csr_mstatus(dcache_io_cpu_tlb_csr_mstatus),
    .io_cpu_tlb_csr_imode(dcache_io_cpu_tlb_csr_imode),
    .io_cpu_tlb_csr_dmode(dcache_io_cpu_tlb_csr_dmode),
    .io_axi_ar_ready(dcache_io_axi_ar_ready),
    .io_axi_ar_valid(dcache_io_axi_ar_valid),
    .io_axi_ar_bits_addr(dcache_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(dcache_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(dcache_io_axi_ar_bits_size),
    .io_axi_r_ready(dcache_io_axi_r_ready),
    .io_axi_r_valid(dcache_io_axi_r_valid),
    .io_axi_r_bits_data(dcache_io_axi_r_bits_data),
    .io_axi_r_bits_resp(dcache_io_axi_r_bits_resp),
    .io_axi_r_bits_last(dcache_io_axi_r_bits_last),
    .io_axi_aw_ready(dcache_io_axi_aw_ready),
    .io_axi_aw_valid(dcache_io_axi_aw_valid),
    .io_axi_aw_bits_addr(dcache_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(dcache_io_axi_aw_bits_len),
    .io_axi_aw_bits_size(dcache_io_axi_aw_bits_size),
    .io_axi_w_ready(dcache_io_axi_w_ready),
    .io_axi_w_valid(dcache_io_axi_w_valid),
    .io_axi_w_bits_data(dcache_io_axi_w_bits_data),
    .io_axi_w_bits_strb(dcache_io_axi_w_bits_strb),
    .io_axi_w_bits_last(dcache_io_axi_w_bits_last),
    .io_axi_b_ready(dcache_io_axi_b_ready),
    .io_axi_b_valid(dcache_io_axi_b_valid)
  );
  CacheAXIInterface axi_interface ( // @[playground/src/cache/Cache.scala 22:29]
    .clock(axi_interface_clock),
    .reset(axi_interface_reset),
    .io_icache_ar_ready(axi_interface_io_icache_ar_ready),
    .io_icache_ar_valid(axi_interface_io_icache_ar_valid),
    .io_icache_ar_bits_addr(axi_interface_io_icache_ar_bits_addr),
    .io_icache_ar_bits_len(axi_interface_io_icache_ar_bits_len),
    .io_icache_ar_bits_size(axi_interface_io_icache_ar_bits_size),
    .io_icache_r_ready(axi_interface_io_icache_r_ready),
    .io_icache_r_valid(axi_interface_io_icache_r_valid),
    .io_icache_r_bits_data(axi_interface_io_icache_r_bits_data),
    .io_icache_r_bits_resp(axi_interface_io_icache_r_bits_resp),
    .io_icache_r_bits_last(axi_interface_io_icache_r_bits_last),
    .io_dcache_ar_ready(axi_interface_io_dcache_ar_ready),
    .io_dcache_ar_valid(axi_interface_io_dcache_ar_valid),
    .io_dcache_ar_bits_addr(axi_interface_io_dcache_ar_bits_addr),
    .io_dcache_ar_bits_len(axi_interface_io_dcache_ar_bits_len),
    .io_dcache_ar_bits_size(axi_interface_io_dcache_ar_bits_size),
    .io_dcache_r_ready(axi_interface_io_dcache_r_ready),
    .io_dcache_r_valid(axi_interface_io_dcache_r_valid),
    .io_dcache_r_bits_data(axi_interface_io_dcache_r_bits_data),
    .io_dcache_r_bits_resp(axi_interface_io_dcache_r_bits_resp),
    .io_dcache_r_bits_last(axi_interface_io_dcache_r_bits_last),
    .io_dcache_aw_ready(axi_interface_io_dcache_aw_ready),
    .io_dcache_aw_valid(axi_interface_io_dcache_aw_valid),
    .io_dcache_aw_bits_addr(axi_interface_io_dcache_aw_bits_addr),
    .io_dcache_aw_bits_len(axi_interface_io_dcache_aw_bits_len),
    .io_dcache_aw_bits_size(axi_interface_io_dcache_aw_bits_size),
    .io_dcache_w_ready(axi_interface_io_dcache_w_ready),
    .io_dcache_w_valid(axi_interface_io_dcache_w_valid),
    .io_dcache_w_bits_data(axi_interface_io_dcache_w_bits_data),
    .io_dcache_w_bits_strb(axi_interface_io_dcache_w_bits_strb),
    .io_dcache_w_bits_last(axi_interface_io_dcache_w_bits_last),
    .io_dcache_b_valid(axi_interface_io_dcache_b_valid),
    .io_axi_ar_ready(axi_interface_io_axi_ar_ready),
    .io_axi_ar_valid(axi_interface_io_axi_ar_valid),
    .io_axi_ar_bits_id(axi_interface_io_axi_ar_bits_id),
    .io_axi_ar_bits_addr(axi_interface_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(axi_interface_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(axi_interface_io_axi_ar_bits_size),
    .io_axi_r_ready(axi_interface_io_axi_r_ready),
    .io_axi_r_valid(axi_interface_io_axi_r_valid),
    .io_axi_r_bits_id(axi_interface_io_axi_r_bits_id),
    .io_axi_r_bits_data(axi_interface_io_axi_r_bits_data),
    .io_axi_r_bits_resp(axi_interface_io_axi_r_bits_resp),
    .io_axi_r_bits_last(axi_interface_io_axi_r_bits_last),
    .io_axi_aw_ready(axi_interface_io_axi_aw_ready),
    .io_axi_aw_valid(axi_interface_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axi_interface_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(axi_interface_io_axi_aw_bits_len),
    .io_axi_aw_bits_size(axi_interface_io_axi_aw_bits_size),
    .io_axi_w_ready(axi_interface_io_axi_w_ready),
    .io_axi_w_valid(axi_interface_io_axi_w_valid),
    .io_axi_w_bits_data(axi_interface_io_axi_w_bits_data),
    .io_axi_w_bits_strb(axi_interface_io_axi_w_bits_strb),
    .io_axi_w_bits_last(axi_interface_io_axi_w_bits_last),
    .io_axi_b_valid(axi_interface_io_axi_b_valid)
  );
  assign io_inst_inst_0 = icache_io_cpu_inst_0; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_inst_1 = icache_io_cpu_inst_1; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_inst_valid_0 = icache_io_cpu_inst_valid_0; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_inst_valid_1 = icache_io_cpu_inst_valid_1; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_access_fault = icache_io_cpu_access_fault; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_page_fault = icache_io_cpu_page_fault; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_addr_misaligned = icache_io_cpu_addr_misaligned; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_icache_stall = icache_io_cpu_icache_stall; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_tlb_en = icache_io_cpu_tlb_en; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_tlb_vaddr = icache_io_cpu_tlb_vaddr; // @[playground/src/cache/Cache.scala 27:11]
  assign io_inst_tlb_complete_single_request = icache_io_cpu_tlb_complete_single_request; // @[playground/src/cache/Cache.scala 27:11]
  assign io_data_rdata = dcache_io_cpu_rdata; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_access_fault = dcache_io_cpu_access_fault; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_page_fault = dcache_io_cpu_page_fault; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_dcache_ready = dcache_io_cpu_dcache_ready; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_en = dcache_io_cpu_tlb_en; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_vaddr = dcache_io_cpu_tlb_vaddr; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_complete_single_request = dcache_io_cpu_tlb_complete_single_request; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_access_type = dcache_io_cpu_tlb_access_type; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_vpn_ready = dcache_io_cpu_tlb_ptw_vpn_ready; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_valid = dcache_io_cpu_tlb_ptw_pte_valid; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_page_fault = dcache_io_cpu_tlb_ptw_pte_bits_page_fault; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_ppn = dcache_io_cpu_tlb_ptw_pte_bits_entry_ppn; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_d = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_d; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_g = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_g; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_u = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_u; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_x = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_x; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_w = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_w; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_r = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_r; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_entry_flag_v = dcache_io_cpu_tlb_ptw_pte_bits_entry_flag_v; // @[playground/src/cache/Cache.scala 28:11]
  assign io_data_tlb_ptw_pte_bits_rmask = dcache_io_cpu_tlb_ptw_pte_bits_rmask; // @[playground/src/cache/Cache.scala 28:11]
  assign io_axi_ar_valid = axi_interface_io_axi_ar_valid; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_ar_bits_id = axi_interface_io_axi_ar_bits_id; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_ar_bits_addr = axi_interface_io_axi_ar_bits_addr; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_ar_bits_len = axi_interface_io_axi_ar_bits_len; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_ar_bits_size = axi_interface_io_axi_ar_bits_size; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_r_ready = axi_interface_io_axi_r_ready; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_aw_valid = axi_interface_io_axi_aw_valid; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_aw_bits_addr = axi_interface_io_axi_aw_bits_addr; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_aw_bits_len = axi_interface_io_axi_aw_bits_len; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_aw_bits_size = axi_interface_io_axi_aw_bits_size; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_w_valid = axi_interface_io_axi_w_valid; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_w_bits_data = axi_interface_io_axi_w_bits_data; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_w_bits_strb = axi_interface_io_axi_w_bits_strb; // @[playground/src/cache/Cache.scala 29:10]
  assign io_axi_w_bits_last = axi_interface_io_axi_w_bits_last; // @[playground/src/cache/Cache.scala 29:10]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_cpu_req = io_inst_req; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_complete_single_request = io_inst_complete_single_request; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_addr_0 = io_inst_addr_0; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_addr_1 = io_inst_addr_1; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_fence_i = io_inst_fence_i; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_dcache_stall = io_inst_dcache_stall; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_tlb_uncached = io_inst_tlb_uncached; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_tlb_hit = io_inst_tlb_hit; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_tlb_ptag = io_inst_tlb_ptag; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_tlb_paddr = io_inst_tlb_paddr; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_cpu_tlb_page_fault = io_inst_tlb_page_fault; // @[playground/src/cache/Cache.scala 27:11]
  assign icache_io_axi_ar_ready = axi_interface_io_icache_ar_ready; // @[playground/src/cache/Cache.scala 24:17]
  assign icache_io_axi_r_valid = axi_interface_io_icache_r_valid; // @[playground/src/cache/Cache.scala 24:17]
  assign icache_io_axi_r_bits_data = axi_interface_io_icache_r_bits_data; // @[playground/src/cache/Cache.scala 24:17]
  assign icache_io_axi_r_bits_resp = axi_interface_io_icache_r_bits_resp; // @[playground/src/cache/Cache.scala 24:17]
  assign icache_io_axi_r_bits_last = axi_interface_io_icache_r_bits_last; // @[playground/src/cache/Cache.scala 24:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_cpu_exe_addr = io_data_exe_addr; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_addr = io_data_addr; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_rlen = io_data_rlen; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_en = io_data_en; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_wen = io_data_wen; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_wdata = io_data_wdata; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_complete_single_request = io_data_complete_single_request; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_fence_i = io_data_fence_i; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_wstrb = io_data_wstrb; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_uncached = io_data_tlb_uncached; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_hit = io_data_tlb_hit; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_ptag = io_data_tlb_ptag; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_paddr = io_data_tlb_paddr; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_page_fault = io_data_tlb_page_fault; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_ptw_vpn_valid = io_data_tlb_ptw_vpn_valid; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_ptw_vpn_bits = io_data_tlb_ptw_vpn_bits; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_ptw_access_type = io_data_tlb_ptw_access_type; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_csr_satp = io_data_tlb_csr_satp; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_csr_mstatus = io_data_tlb_csr_mstatus; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_csr_imode = io_data_tlb_csr_imode; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_cpu_tlb_csr_dmode = io_data_tlb_csr_dmode; // @[playground/src/cache/Cache.scala 28:11]
  assign dcache_io_axi_ar_ready = axi_interface_io_dcache_ar_ready; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_r_valid = axi_interface_io_dcache_r_valid; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_r_bits_data = axi_interface_io_dcache_r_bits_data; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_r_bits_resp = axi_interface_io_dcache_r_bits_resp; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_r_bits_last = axi_interface_io_dcache_r_bits_last; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_aw_ready = axi_interface_io_dcache_aw_ready; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_w_ready = axi_interface_io_dcache_w_ready; // @[playground/src/cache/Cache.scala 25:17]
  assign dcache_io_axi_b_valid = axi_interface_io_dcache_b_valid; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_clock = clock;
  assign axi_interface_reset = reset;
  assign axi_interface_io_icache_ar_valid = icache_io_axi_ar_valid; // @[playground/src/cache/Cache.scala 24:17]
  assign axi_interface_io_icache_ar_bits_addr = icache_io_axi_ar_bits_addr; // @[playground/src/cache/Cache.scala 24:17]
  assign axi_interface_io_icache_ar_bits_len = icache_io_axi_ar_bits_len; // @[playground/src/cache/Cache.scala 24:17]
  assign axi_interface_io_icache_ar_bits_size = icache_io_axi_ar_bits_size; // @[playground/src/cache/Cache.scala 24:17]
  assign axi_interface_io_icache_r_ready = icache_io_axi_r_ready; // @[playground/src/cache/Cache.scala 24:17]
  assign axi_interface_io_dcache_ar_valid = dcache_io_axi_ar_valid; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_ar_bits_addr = dcache_io_axi_ar_bits_addr; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_ar_bits_len = dcache_io_axi_ar_bits_len; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_ar_bits_size = dcache_io_axi_ar_bits_size; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_r_ready = dcache_io_axi_r_ready; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_aw_valid = dcache_io_axi_aw_valid; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_aw_bits_addr = dcache_io_axi_aw_bits_addr; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_aw_bits_len = dcache_io_axi_aw_bits_len; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_aw_bits_size = dcache_io_axi_aw_bits_size; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_w_valid = dcache_io_axi_w_valid; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_w_bits_data = dcache_io_axi_w_bits_data; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_w_bits_strb = dcache_io_axi_w_bits_strb; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_dcache_w_bits_last = dcache_io_axi_w_bits_last; // @[playground/src/cache/Cache.scala 25:17]
  assign axi_interface_io_axi_ar_ready = io_axi_ar_ready; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_r_valid = io_axi_r_valid; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_r_bits_id = io_axi_r_bits_id; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_r_bits_data = io_axi_r_bits_data; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_r_bits_resp = io_axi_r_bits_resp; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_r_bits_last = io_axi_r_bits_last; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_aw_ready = io_axi_aw_ready; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_w_ready = io_axi_w_ready; // @[playground/src/cache/Cache.scala 29:10]
  assign axi_interface_io_axi_b_valid = io_axi_b_valid; // @[playground/src/cache/Cache.scala 29:10]
endmodule
module PuaCpu(
  input         clock,
  input         reset,
  input         io_ext_int_ei, // @[playground/src/PuaCpu.scala 9:14]
  input         io_ext_int_ti, // @[playground/src/PuaCpu.scala 9:14]
  input         io_ext_int_si, // @[playground/src/PuaCpu.scala 9:14]
  input         io_axi_ar_ready, // @[playground/src/PuaCpu.scala 9:14]
  output        io_axi_ar_valid, // @[playground/src/PuaCpu.scala 9:14]
  output [3:0]  io_axi_ar_bits_id, // @[playground/src/PuaCpu.scala 9:14]
  output [31:0] io_axi_ar_bits_addr, // @[playground/src/PuaCpu.scala 9:14]
  output [7:0]  io_axi_ar_bits_len, // @[playground/src/PuaCpu.scala 9:14]
  output [2:0]  io_axi_ar_bits_size, // @[playground/src/PuaCpu.scala 9:14]
  output [1:0]  io_axi_ar_bits_burst, // @[playground/src/PuaCpu.scala 9:14]
  output [1:0]  io_axi_ar_bits_lock, // @[playground/src/PuaCpu.scala 9:14]
  output [3:0]  io_axi_ar_bits_cache, // @[playground/src/PuaCpu.scala 9:14]
  output [2:0]  io_axi_ar_bits_prot, // @[playground/src/PuaCpu.scala 9:14]
  output        io_axi_r_ready, // @[playground/src/PuaCpu.scala 9:14]
  input         io_axi_r_valid, // @[playground/src/PuaCpu.scala 9:14]
  input  [3:0]  io_axi_r_bits_id, // @[playground/src/PuaCpu.scala 9:14]
  input  [63:0] io_axi_r_bits_data, // @[playground/src/PuaCpu.scala 9:14]
  input  [1:0]  io_axi_r_bits_resp, // @[playground/src/PuaCpu.scala 9:14]
  input         io_axi_r_bits_last, // @[playground/src/PuaCpu.scala 9:14]
  input         io_axi_aw_ready, // @[playground/src/PuaCpu.scala 9:14]
  output        io_axi_aw_valid, // @[playground/src/PuaCpu.scala 9:14]
  output [3:0]  io_axi_aw_bits_id, // @[playground/src/PuaCpu.scala 9:14]
  output [31:0] io_axi_aw_bits_addr, // @[playground/src/PuaCpu.scala 9:14]
  output [7:0]  io_axi_aw_bits_len, // @[playground/src/PuaCpu.scala 9:14]
  output [2:0]  io_axi_aw_bits_size, // @[playground/src/PuaCpu.scala 9:14]
  output [1:0]  io_axi_aw_bits_burst, // @[playground/src/PuaCpu.scala 9:14]
  output [1:0]  io_axi_aw_bits_lock, // @[playground/src/PuaCpu.scala 9:14]
  output [3:0]  io_axi_aw_bits_cache, // @[playground/src/PuaCpu.scala 9:14]
  output [2:0]  io_axi_aw_bits_prot, // @[playground/src/PuaCpu.scala 9:14]
  input         io_axi_w_ready, // @[playground/src/PuaCpu.scala 9:14]
  output        io_axi_w_valid, // @[playground/src/PuaCpu.scala 9:14]
  output [3:0]  io_axi_w_bits_id, // @[playground/src/PuaCpu.scala 9:14]
  output [63:0] io_axi_w_bits_data, // @[playground/src/PuaCpu.scala 9:14]
  output [7:0]  io_axi_w_bits_strb, // @[playground/src/PuaCpu.scala 9:14]
  output        io_axi_w_bits_last, // @[playground/src/PuaCpu.scala 9:14]
  output        io_axi_b_ready, // @[playground/src/PuaCpu.scala 9:14]
  input         io_axi_b_valid, // @[playground/src/PuaCpu.scala 9:14]
  input  [3:0]  io_axi_b_bits_id, // @[playground/src/PuaCpu.scala 9:14]
  input  [1:0]  io_axi_b_bits_resp, // @[playground/src/PuaCpu.scala 9:14]
  output [63:0] io_debug_wb_pc, // @[playground/src/PuaCpu.scala 9:14]
  output        io_debug_wb_rf_wen, // @[playground/src/PuaCpu.scala 9:14]
  output [4:0]  io_debug_wb_rf_wnum, // @[playground/src/PuaCpu.scala 9:14]
  output [63:0] io_debug_wb_rf_wdata // @[playground/src/PuaCpu.scala 9:14]
);
  wire  core_clock; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_reset; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_ext_int_ei; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_ext_int_ti; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_ext_int_si; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_req; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_complete_single_request; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_inst_addr_0; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_inst_addr_1; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_fence_i; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_dcache_stall; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_inst_inst_0; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_inst_inst_1; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_inst_valid_0; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_inst_valid_1; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_access_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_page_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_addr_misaligned; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_icache_stall; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_tlb_en; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_inst_tlb_vaddr; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_tlb_complete_single_request; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_tlb_uncached; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_tlb_hit; // @[playground/src/PuaCpu.scala 14:21]
  wire [19:0] core_io_inst_tlb_ptag; // @[playground/src/PuaCpu.scala 14:21]
  wire [31:0] core_io_inst_tlb_paddr; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_inst_tlb_page_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_exe_addr; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_addr; // @[playground/src/PuaCpu.scala 14:21]
  wire [7:0] core_io_data_rlen; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_en; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_wen; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_wdata; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_complete_single_request; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_fence_i; // @[playground/src/PuaCpu.scala 14:21]
  wire [7:0] core_io_data_wstrb; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_rdata; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_access_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_page_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_dcache_ready; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_en; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_tlb_vaddr; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_complete_single_request; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_uncached; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_hit; // @[playground/src/PuaCpu.scala 14:21]
  wire [19:0] core_io_data_tlb_ptag; // @[playground/src/PuaCpu.scala 14:21]
  wire [31:0] core_io_data_tlb_paddr; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_page_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire [1:0] core_io_data_tlb_access_type; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_vpn_ready; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_vpn_valid; // @[playground/src/PuaCpu.scala 14:21]
  wire [26:0] core_io_data_tlb_ptw_vpn_bits; // @[playground/src/PuaCpu.scala 14:21]
  wire [1:0] core_io_data_tlb_ptw_access_type; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_valid; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_page_fault; // @[playground/src/PuaCpu.scala 14:21]
  wire [19:0] core_io_data_tlb_ptw_pte_bits_entry_ppn; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_d; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_g; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_u; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_x; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_w; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_r; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_data_tlb_ptw_pte_bits_entry_flag_v; // @[playground/src/PuaCpu.scala 14:21]
  wire [17:0] core_io_data_tlb_ptw_pte_bits_rmask; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_tlb_csr_satp; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_data_tlb_csr_mstatus; // @[playground/src/PuaCpu.scala 14:21]
  wire [1:0] core_io_data_tlb_csr_imode; // @[playground/src/PuaCpu.scala 14:21]
  wire [1:0] core_io_data_tlb_csr_dmode; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_debug_wb_pc; // @[playground/src/PuaCpu.scala 14:21]
  wire  core_io_debug_wb_rf_wen; // @[playground/src/PuaCpu.scala 14:21]
  wire [4:0] core_io_debug_wb_rf_wnum; // @[playground/src/PuaCpu.scala 14:21]
  wire [63:0] core_io_debug_wb_rf_wdata; // @[playground/src/PuaCpu.scala 14:21]
  wire  cache_clock; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_reset; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_req; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_complete_single_request; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_inst_addr_0; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_inst_addr_1; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_fence_i; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_dcache_stall; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_inst_inst_0; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_inst_inst_1; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_inst_valid_0; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_inst_valid_1; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_access_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_page_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_addr_misaligned; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_icache_stall; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_tlb_en; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_inst_tlb_vaddr; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_tlb_complete_single_request; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_tlb_uncached; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_tlb_hit; // @[playground/src/PuaCpu.scala 15:21]
  wire [19:0] cache_io_inst_tlb_ptag; // @[playground/src/PuaCpu.scala 15:21]
  wire [31:0] cache_io_inst_tlb_paddr; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_inst_tlb_page_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_exe_addr; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_addr; // @[playground/src/PuaCpu.scala 15:21]
  wire [7:0] cache_io_data_rlen; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_en; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_wen; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_wdata; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_complete_single_request; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_fence_i; // @[playground/src/PuaCpu.scala 15:21]
  wire [7:0] cache_io_data_wstrb; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_rdata; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_access_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_page_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_dcache_ready; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_en; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_tlb_vaddr; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_complete_single_request; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_uncached; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_hit; // @[playground/src/PuaCpu.scala 15:21]
  wire [19:0] cache_io_data_tlb_ptag; // @[playground/src/PuaCpu.scala 15:21]
  wire [31:0] cache_io_data_tlb_paddr; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_page_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire [1:0] cache_io_data_tlb_access_type; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_vpn_ready; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_vpn_valid; // @[playground/src/PuaCpu.scala 15:21]
  wire [26:0] cache_io_data_tlb_ptw_vpn_bits; // @[playground/src/PuaCpu.scala 15:21]
  wire [1:0] cache_io_data_tlb_ptw_access_type; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_valid; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_page_fault; // @[playground/src/PuaCpu.scala 15:21]
  wire [19:0] cache_io_data_tlb_ptw_pte_bits_entry_ppn; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_d; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_g; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_u; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_x; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_w; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_r; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_data_tlb_ptw_pte_bits_entry_flag_v; // @[playground/src/PuaCpu.scala 15:21]
  wire [17:0] cache_io_data_tlb_ptw_pte_bits_rmask; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_tlb_csr_satp; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_data_tlb_csr_mstatus; // @[playground/src/PuaCpu.scala 15:21]
  wire [1:0] cache_io_data_tlb_csr_imode; // @[playground/src/PuaCpu.scala 15:21]
  wire [1:0] cache_io_data_tlb_csr_dmode; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_ar_ready; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_ar_valid; // @[playground/src/PuaCpu.scala 15:21]
  wire [3:0] cache_io_axi_ar_bits_id; // @[playground/src/PuaCpu.scala 15:21]
  wire [31:0] cache_io_axi_ar_bits_addr; // @[playground/src/PuaCpu.scala 15:21]
  wire [7:0] cache_io_axi_ar_bits_len; // @[playground/src/PuaCpu.scala 15:21]
  wire [2:0] cache_io_axi_ar_bits_size; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_r_ready; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_r_valid; // @[playground/src/PuaCpu.scala 15:21]
  wire [3:0] cache_io_axi_r_bits_id; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_axi_r_bits_data; // @[playground/src/PuaCpu.scala 15:21]
  wire [1:0] cache_io_axi_r_bits_resp; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_r_bits_last; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_aw_ready; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_aw_valid; // @[playground/src/PuaCpu.scala 15:21]
  wire [31:0] cache_io_axi_aw_bits_addr; // @[playground/src/PuaCpu.scala 15:21]
  wire [7:0] cache_io_axi_aw_bits_len; // @[playground/src/PuaCpu.scala 15:21]
  wire [2:0] cache_io_axi_aw_bits_size; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_w_ready; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_w_valid; // @[playground/src/PuaCpu.scala 15:21]
  wire [63:0] cache_io_axi_w_bits_data; // @[playground/src/PuaCpu.scala 15:21]
  wire [7:0] cache_io_axi_w_bits_strb; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_w_bits_last; // @[playground/src/PuaCpu.scala 15:21]
  wire  cache_io_axi_b_valid; // @[playground/src/PuaCpu.scala 15:21]
  Core core ( // @[playground/src/PuaCpu.scala 14:21]
    .clock(core_clock),
    .reset(core_reset),
    .io_ext_int_ei(core_io_ext_int_ei),
    .io_ext_int_ti(core_io_ext_int_ti),
    .io_ext_int_si(core_io_ext_int_si),
    .io_inst_req(core_io_inst_req),
    .io_inst_complete_single_request(core_io_inst_complete_single_request),
    .io_inst_addr_0(core_io_inst_addr_0),
    .io_inst_addr_1(core_io_inst_addr_1),
    .io_inst_fence_i(core_io_inst_fence_i),
    .io_inst_dcache_stall(core_io_inst_dcache_stall),
    .io_inst_inst_0(core_io_inst_inst_0),
    .io_inst_inst_1(core_io_inst_inst_1),
    .io_inst_inst_valid_0(core_io_inst_inst_valid_0),
    .io_inst_inst_valid_1(core_io_inst_inst_valid_1),
    .io_inst_access_fault(core_io_inst_access_fault),
    .io_inst_page_fault(core_io_inst_page_fault),
    .io_inst_addr_misaligned(core_io_inst_addr_misaligned),
    .io_inst_icache_stall(core_io_inst_icache_stall),
    .io_inst_tlb_en(core_io_inst_tlb_en),
    .io_inst_tlb_vaddr(core_io_inst_tlb_vaddr),
    .io_inst_tlb_complete_single_request(core_io_inst_tlb_complete_single_request),
    .io_inst_tlb_uncached(core_io_inst_tlb_uncached),
    .io_inst_tlb_hit(core_io_inst_tlb_hit),
    .io_inst_tlb_ptag(core_io_inst_tlb_ptag),
    .io_inst_tlb_paddr(core_io_inst_tlb_paddr),
    .io_inst_tlb_page_fault(core_io_inst_tlb_page_fault),
    .io_data_exe_addr(core_io_data_exe_addr),
    .io_data_addr(core_io_data_addr),
    .io_data_rlen(core_io_data_rlen),
    .io_data_en(core_io_data_en),
    .io_data_wen(core_io_data_wen),
    .io_data_wdata(core_io_data_wdata),
    .io_data_complete_single_request(core_io_data_complete_single_request),
    .io_data_fence_i(core_io_data_fence_i),
    .io_data_wstrb(core_io_data_wstrb),
    .io_data_rdata(core_io_data_rdata),
    .io_data_access_fault(core_io_data_access_fault),
    .io_data_page_fault(core_io_data_page_fault),
    .io_data_dcache_ready(core_io_data_dcache_ready),
    .io_data_tlb_en(core_io_data_tlb_en),
    .io_data_tlb_vaddr(core_io_data_tlb_vaddr),
    .io_data_tlb_complete_single_request(core_io_data_tlb_complete_single_request),
    .io_data_tlb_uncached(core_io_data_tlb_uncached),
    .io_data_tlb_hit(core_io_data_tlb_hit),
    .io_data_tlb_ptag(core_io_data_tlb_ptag),
    .io_data_tlb_paddr(core_io_data_tlb_paddr),
    .io_data_tlb_page_fault(core_io_data_tlb_page_fault),
    .io_data_tlb_access_type(core_io_data_tlb_access_type),
    .io_data_tlb_ptw_vpn_ready(core_io_data_tlb_ptw_vpn_ready),
    .io_data_tlb_ptw_vpn_valid(core_io_data_tlb_ptw_vpn_valid),
    .io_data_tlb_ptw_vpn_bits(core_io_data_tlb_ptw_vpn_bits),
    .io_data_tlb_ptw_access_type(core_io_data_tlb_ptw_access_type),
    .io_data_tlb_ptw_pte_valid(core_io_data_tlb_ptw_pte_valid),
    .io_data_tlb_ptw_pte_bits_page_fault(core_io_data_tlb_ptw_pte_bits_page_fault),
    .io_data_tlb_ptw_pte_bits_entry_ppn(core_io_data_tlb_ptw_pte_bits_entry_ppn),
    .io_data_tlb_ptw_pte_bits_entry_flag_d(core_io_data_tlb_ptw_pte_bits_entry_flag_d),
    .io_data_tlb_ptw_pte_bits_entry_flag_g(core_io_data_tlb_ptw_pte_bits_entry_flag_g),
    .io_data_tlb_ptw_pte_bits_entry_flag_u(core_io_data_tlb_ptw_pte_bits_entry_flag_u),
    .io_data_tlb_ptw_pte_bits_entry_flag_x(core_io_data_tlb_ptw_pte_bits_entry_flag_x),
    .io_data_tlb_ptw_pte_bits_entry_flag_w(core_io_data_tlb_ptw_pte_bits_entry_flag_w),
    .io_data_tlb_ptw_pte_bits_entry_flag_r(core_io_data_tlb_ptw_pte_bits_entry_flag_r),
    .io_data_tlb_ptw_pte_bits_entry_flag_v(core_io_data_tlb_ptw_pte_bits_entry_flag_v),
    .io_data_tlb_ptw_pte_bits_rmask(core_io_data_tlb_ptw_pte_bits_rmask),
    .io_data_tlb_csr_satp(core_io_data_tlb_csr_satp),
    .io_data_tlb_csr_mstatus(core_io_data_tlb_csr_mstatus),
    .io_data_tlb_csr_imode(core_io_data_tlb_csr_imode),
    .io_data_tlb_csr_dmode(core_io_data_tlb_csr_dmode),
    .io_debug_wb_pc(core_io_debug_wb_pc),
    .io_debug_wb_rf_wen(core_io_debug_wb_rf_wen),
    .io_debug_wb_rf_wnum(core_io_debug_wb_rf_wnum),
    .io_debug_wb_rf_wdata(core_io_debug_wb_rf_wdata)
  );
  Cache cache ( // @[playground/src/PuaCpu.scala 15:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_inst_req(cache_io_inst_req),
    .io_inst_complete_single_request(cache_io_inst_complete_single_request),
    .io_inst_addr_0(cache_io_inst_addr_0),
    .io_inst_addr_1(cache_io_inst_addr_1),
    .io_inst_fence_i(cache_io_inst_fence_i),
    .io_inst_dcache_stall(cache_io_inst_dcache_stall),
    .io_inst_inst_0(cache_io_inst_inst_0),
    .io_inst_inst_1(cache_io_inst_inst_1),
    .io_inst_inst_valid_0(cache_io_inst_inst_valid_0),
    .io_inst_inst_valid_1(cache_io_inst_inst_valid_1),
    .io_inst_access_fault(cache_io_inst_access_fault),
    .io_inst_page_fault(cache_io_inst_page_fault),
    .io_inst_addr_misaligned(cache_io_inst_addr_misaligned),
    .io_inst_icache_stall(cache_io_inst_icache_stall),
    .io_inst_tlb_en(cache_io_inst_tlb_en),
    .io_inst_tlb_vaddr(cache_io_inst_tlb_vaddr),
    .io_inst_tlb_complete_single_request(cache_io_inst_tlb_complete_single_request),
    .io_inst_tlb_uncached(cache_io_inst_tlb_uncached),
    .io_inst_tlb_hit(cache_io_inst_tlb_hit),
    .io_inst_tlb_ptag(cache_io_inst_tlb_ptag),
    .io_inst_tlb_paddr(cache_io_inst_tlb_paddr),
    .io_inst_tlb_page_fault(cache_io_inst_tlb_page_fault),
    .io_data_exe_addr(cache_io_data_exe_addr),
    .io_data_addr(cache_io_data_addr),
    .io_data_rlen(cache_io_data_rlen),
    .io_data_en(cache_io_data_en),
    .io_data_wen(cache_io_data_wen),
    .io_data_wdata(cache_io_data_wdata),
    .io_data_complete_single_request(cache_io_data_complete_single_request),
    .io_data_fence_i(cache_io_data_fence_i),
    .io_data_wstrb(cache_io_data_wstrb),
    .io_data_rdata(cache_io_data_rdata),
    .io_data_access_fault(cache_io_data_access_fault),
    .io_data_page_fault(cache_io_data_page_fault),
    .io_data_dcache_ready(cache_io_data_dcache_ready),
    .io_data_tlb_en(cache_io_data_tlb_en),
    .io_data_tlb_vaddr(cache_io_data_tlb_vaddr),
    .io_data_tlb_complete_single_request(cache_io_data_tlb_complete_single_request),
    .io_data_tlb_uncached(cache_io_data_tlb_uncached),
    .io_data_tlb_hit(cache_io_data_tlb_hit),
    .io_data_tlb_ptag(cache_io_data_tlb_ptag),
    .io_data_tlb_paddr(cache_io_data_tlb_paddr),
    .io_data_tlb_page_fault(cache_io_data_tlb_page_fault),
    .io_data_tlb_access_type(cache_io_data_tlb_access_type),
    .io_data_tlb_ptw_vpn_ready(cache_io_data_tlb_ptw_vpn_ready),
    .io_data_tlb_ptw_vpn_valid(cache_io_data_tlb_ptw_vpn_valid),
    .io_data_tlb_ptw_vpn_bits(cache_io_data_tlb_ptw_vpn_bits),
    .io_data_tlb_ptw_access_type(cache_io_data_tlb_ptw_access_type),
    .io_data_tlb_ptw_pte_valid(cache_io_data_tlb_ptw_pte_valid),
    .io_data_tlb_ptw_pte_bits_page_fault(cache_io_data_tlb_ptw_pte_bits_page_fault),
    .io_data_tlb_ptw_pte_bits_entry_ppn(cache_io_data_tlb_ptw_pte_bits_entry_ppn),
    .io_data_tlb_ptw_pte_bits_entry_flag_d(cache_io_data_tlb_ptw_pte_bits_entry_flag_d),
    .io_data_tlb_ptw_pte_bits_entry_flag_g(cache_io_data_tlb_ptw_pte_bits_entry_flag_g),
    .io_data_tlb_ptw_pte_bits_entry_flag_u(cache_io_data_tlb_ptw_pte_bits_entry_flag_u),
    .io_data_tlb_ptw_pte_bits_entry_flag_x(cache_io_data_tlb_ptw_pte_bits_entry_flag_x),
    .io_data_tlb_ptw_pte_bits_entry_flag_w(cache_io_data_tlb_ptw_pte_bits_entry_flag_w),
    .io_data_tlb_ptw_pte_bits_entry_flag_r(cache_io_data_tlb_ptw_pte_bits_entry_flag_r),
    .io_data_tlb_ptw_pte_bits_entry_flag_v(cache_io_data_tlb_ptw_pte_bits_entry_flag_v),
    .io_data_tlb_ptw_pte_bits_rmask(cache_io_data_tlb_ptw_pte_bits_rmask),
    .io_data_tlb_csr_satp(cache_io_data_tlb_csr_satp),
    .io_data_tlb_csr_mstatus(cache_io_data_tlb_csr_mstatus),
    .io_data_tlb_csr_imode(cache_io_data_tlb_csr_imode),
    .io_data_tlb_csr_dmode(cache_io_data_tlb_csr_dmode),
    .io_axi_ar_ready(cache_io_axi_ar_ready),
    .io_axi_ar_valid(cache_io_axi_ar_valid),
    .io_axi_ar_bits_id(cache_io_axi_ar_bits_id),
    .io_axi_ar_bits_addr(cache_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(cache_io_axi_ar_bits_len),
    .io_axi_ar_bits_size(cache_io_axi_ar_bits_size),
    .io_axi_r_ready(cache_io_axi_r_ready),
    .io_axi_r_valid(cache_io_axi_r_valid),
    .io_axi_r_bits_id(cache_io_axi_r_bits_id),
    .io_axi_r_bits_data(cache_io_axi_r_bits_data),
    .io_axi_r_bits_resp(cache_io_axi_r_bits_resp),
    .io_axi_r_bits_last(cache_io_axi_r_bits_last),
    .io_axi_aw_ready(cache_io_axi_aw_ready),
    .io_axi_aw_valid(cache_io_axi_aw_valid),
    .io_axi_aw_bits_addr(cache_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(cache_io_axi_aw_bits_len),
    .io_axi_aw_bits_size(cache_io_axi_aw_bits_size),
    .io_axi_w_ready(cache_io_axi_w_ready),
    .io_axi_w_valid(cache_io_axi_w_valid),
    .io_axi_w_bits_data(cache_io_axi_w_bits_data),
    .io_axi_w_bits_strb(cache_io_axi_w_bits_strb),
    .io_axi_w_bits_last(cache_io_axi_w_bits_last),
    .io_axi_b_valid(cache_io_axi_b_valid)
  );
  assign io_axi_ar_valid = cache_io_axi_ar_valid; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_id = cache_io_axi_ar_bits_id; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_addr = cache_io_axi_ar_bits_addr; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_len = cache_io_axi_ar_bits_len; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_size = cache_io_axi_ar_bits_size; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_burst = 2'h1; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_lock = 2'h0; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_cache = 4'h0; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_ar_bits_prot = 3'h0; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_r_ready = cache_io_axi_r_ready; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_valid = cache_io_axi_aw_valid; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_id = 4'h1; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_addr = cache_io_axi_aw_bits_addr; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_len = cache_io_axi_aw_bits_len; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_size = cache_io_axi_aw_bits_size; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_burst = 2'h1; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_lock = 2'h0; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_cache = 4'h0; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_aw_bits_prot = 3'h0; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_w_valid = cache_io_axi_w_valid; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_w_bits_id = 4'h1; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_w_bits_data = cache_io_axi_w_bits_data; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_w_bits_strb = cache_io_axi_w_bits_strb; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_w_bits_last = cache_io_axi_w_bits_last; // @[playground/src/PuaCpu.scala 22:10]
  assign io_axi_b_ready = 1'h1; // @[playground/src/PuaCpu.scala 22:10]
  assign io_debug_wb_pc = core_io_debug_wb_pc; // @[playground/src/PuaCpu.scala 21:12]
  assign io_debug_wb_rf_wen = core_io_debug_wb_rf_wen; // @[playground/src/PuaCpu.scala 21:12]
  assign io_debug_wb_rf_wnum = core_io_debug_wb_rf_wnum; // @[playground/src/PuaCpu.scala 21:12]
  assign io_debug_wb_rf_wdata = core_io_debug_wb_rf_wdata; // @[playground/src/PuaCpu.scala 21:12]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_ext_int_ei = io_ext_int_ei; // @[playground/src/PuaCpu.scala 20:14]
  assign core_io_ext_int_ti = io_ext_int_ti; // @[playground/src/PuaCpu.scala 20:14]
  assign core_io_ext_int_si = io_ext_int_si; // @[playground/src/PuaCpu.scala 20:14]
  assign core_io_inst_inst_0 = cache_io_inst_inst_0; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_inst_1 = cache_io_inst_inst_1; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_inst_valid_0 = cache_io_inst_inst_valid_0; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_inst_valid_1 = cache_io_inst_inst_valid_1; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_access_fault = cache_io_inst_access_fault; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_page_fault = cache_io_inst_page_fault; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_addr_misaligned = cache_io_inst_addr_misaligned; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_icache_stall = cache_io_inst_icache_stall; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_tlb_en = cache_io_inst_tlb_en; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_tlb_vaddr = cache_io_inst_tlb_vaddr; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_inst_tlb_complete_single_request = cache_io_inst_tlb_complete_single_request; // @[playground/src/PuaCpu.scala 17:16]
  assign core_io_data_rdata = cache_io_data_rdata; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_access_fault = cache_io_data_access_fault; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_page_fault = cache_io_data_page_fault; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_dcache_ready = cache_io_data_dcache_ready; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_en = cache_io_data_tlb_en; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_vaddr = cache_io_data_tlb_vaddr; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_complete_single_request = cache_io_data_tlb_complete_single_request; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_access_type = cache_io_data_tlb_access_type; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_vpn_ready = cache_io_data_tlb_ptw_vpn_ready; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_valid = cache_io_data_tlb_ptw_pte_valid; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_page_fault = cache_io_data_tlb_ptw_pte_bits_page_fault; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_ppn = cache_io_data_tlb_ptw_pte_bits_entry_ppn; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_d = cache_io_data_tlb_ptw_pte_bits_entry_flag_d; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_g = cache_io_data_tlb_ptw_pte_bits_entry_flag_g; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_u = cache_io_data_tlb_ptw_pte_bits_entry_flag_u; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_x = cache_io_data_tlb_ptw_pte_bits_entry_flag_x; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_w = cache_io_data_tlb_ptw_pte_bits_entry_flag_w; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_r = cache_io_data_tlb_ptw_pte_bits_entry_flag_r; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_entry_flag_v = cache_io_data_tlb_ptw_pte_bits_entry_flag_v; // @[playground/src/PuaCpu.scala 18:16]
  assign core_io_data_tlb_ptw_pte_bits_rmask = cache_io_data_tlb_ptw_pte_bits_rmask; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_inst_req = core_io_inst_req; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_complete_single_request = core_io_inst_complete_single_request; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_addr_0 = core_io_inst_addr_0; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_addr_1 = core_io_inst_addr_1; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_fence_i = core_io_inst_fence_i; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_dcache_stall = core_io_inst_dcache_stall; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_tlb_uncached = core_io_inst_tlb_uncached; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_tlb_hit = core_io_inst_tlb_hit; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_tlb_ptag = core_io_inst_tlb_ptag; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_tlb_paddr = core_io_inst_tlb_paddr; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_inst_tlb_page_fault = core_io_inst_tlb_page_fault; // @[playground/src/PuaCpu.scala 17:16]
  assign cache_io_data_exe_addr = core_io_data_exe_addr; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_addr = core_io_data_addr; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_rlen = core_io_data_rlen; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_en = core_io_data_en; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_wen = core_io_data_wen; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_wdata = core_io_data_wdata; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_complete_single_request = core_io_data_complete_single_request; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_fence_i = core_io_data_fence_i; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_wstrb = core_io_data_wstrb; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_uncached = core_io_data_tlb_uncached; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_hit = core_io_data_tlb_hit; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_ptag = core_io_data_tlb_ptag; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_paddr = core_io_data_tlb_paddr; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_page_fault = core_io_data_tlb_page_fault; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_ptw_vpn_valid = core_io_data_tlb_ptw_vpn_valid; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_ptw_vpn_bits = core_io_data_tlb_ptw_vpn_bits; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_ptw_access_type = core_io_data_tlb_ptw_access_type; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_csr_satp = core_io_data_tlb_csr_satp; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_csr_mstatus = core_io_data_tlb_csr_mstatus; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_csr_imode = core_io_data_tlb_csr_imode; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_data_tlb_csr_dmode = core_io_data_tlb_csr_dmode; // @[playground/src/PuaCpu.scala 18:16]
  assign cache_io_axi_ar_ready = io_axi_ar_ready; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_r_valid = io_axi_r_valid; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_r_bits_id = io_axi_r_bits_id; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_r_bits_data = io_axi_r_bits_data; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_r_bits_resp = io_axi_r_bits_resp; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_r_bits_last = io_axi_r_bits_last; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_aw_ready = io_axi_aw_ready; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_w_ready = io_axi_w_ready; // @[playground/src/PuaCpu.scala 22:10]
  assign cache_io_axi_b_valid = io_axi_b_valid; // @[playground/src/PuaCpu.scala 22:10]
endmodule
